//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9.03 Education (64-bit)
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Device Version: C
//Created Time: Sun Sep 22 18:32:43 2024

module cart_prom (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [14:0] ad;

wire lut_f_0;
wire lut_f_1;
wire [30:0] prom_inst_0_dout_w;
wire [0:0] prom_inst_0_dout;
wire [30:0] prom_inst_1_dout_w;
wire [0:0] prom_inst_1_dout;
wire [30:0] prom_inst_2_dout_w;
wire [1:1] prom_inst_2_dout;
wire [30:0] prom_inst_3_dout_w;
wire [1:1] prom_inst_3_dout;
wire [30:0] prom_inst_4_dout_w;
wire [2:2] prom_inst_4_dout;
wire [30:0] prom_inst_5_dout_w;
wire [2:2] prom_inst_5_dout;
wire [30:0] prom_inst_6_dout_w;
wire [3:3] prom_inst_6_dout;
wire [30:0] prom_inst_7_dout_w;
wire [3:3] prom_inst_7_dout;
wire [30:0] prom_inst_8_dout_w;
wire [4:4] prom_inst_8_dout;
wire [30:0] prom_inst_9_dout_w;
wire [4:4] prom_inst_9_dout;
wire [30:0] prom_inst_10_dout_w;
wire [5:5] prom_inst_10_dout;
wire [30:0] prom_inst_11_dout_w;
wire [5:5] prom_inst_11_dout;
wire [30:0] prom_inst_12_dout_w;
wire [6:6] prom_inst_12_dout;
wire [30:0] prom_inst_13_dout_w;
wire [6:6] prom_inst_13_dout;
wire [30:0] prom_inst_14_dout_w;
wire [7:7] prom_inst_14_dout;
wire [30:0] prom_inst_15_dout_w;
wire [7:7] prom_inst_15_dout;
wire dff_q_0;

LUT2 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[14])
);
defparam lut_inst_0.INIT = 4'h2;
LUT2 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[14])
);
defparam lut_inst_1.INIT = 4'h8;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],prom_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hFFFFFFFFFFA281D28A154A294D22A2B00A8137C9FBF9F9FDFFFEA7FFFFFFF901;
defparam prom_inst_0.INIT_RAM_01 = 256'hA8B64D9041ACB2CB3EFBEFB7DB5A2513F216116142B998000327D0FF02C8BA2A;
defparam prom_inst_0.INIT_RAM_02 = 256'h1636D46AD15514D22C220ABF21811487489E90723F8A42C104001446B520FFC2;
defparam prom_inst_0.INIT_RAM_03 = 256'h006FE40D96C08F6EAA0A7086D02680810DBDF35FDF6F95FB1CC38CE8F9F48352;
defparam prom_inst_0.INIT_RAM_04 = 256'h80D10CC20C1A85450048C8DA2620512B49A95EF98220A0A2000822914900A8A4;
defparam prom_inst_0.INIT_RAM_05 = 256'h856BD1054607550D8324130C0A694526B20B182454C1A2930200B82AB8294A96;
defparam prom_inst_0.INIT_RAM_06 = 256'h88ACD19E725F420251054BD79E69D1B7554D8C5954450CE942C1450A3774F964;
defparam prom_inst_0.INIT_RAM_07 = 256'h002AA9B32AAAA44456906200DB422B6D0AA0942241C7A4D01052A9888008801A;
defparam prom_inst_0.INIT_RAM_08 = 256'h512655844004400D51170C98C1A2681CB259E374FD5B6D6E822A013E5DEB0000;
defparam prom_inst_0.INIT_RAM_09 = 256'hA6A62256D5511442A1412650A2252A854492540B7EFB200924D1768509284AA1;
defparam prom_inst_0.INIT_RAM_0A = 256'h07960A2385AB914ACC00728791901B1502090A811A5540A24CAA0440D540A24D;
defparam prom_inst_0.INIT_RAM_0B = 256'h0494B8D5A2B01078B17BD8844CD0A20D515155151BBF4B2C413528A24D64902B;
defparam prom_inst_0.INIT_RAM_0C = 256'h0555269073303BE799044E9E64276028A0AAA0AA2A82D2AA88C52C94C455DC54;
defparam prom_inst_0.INIT_RAM_0D = 256'h4088615D658074B692AEF0541510704AB254A1C1B158FA9F9592414057C10050;
defparam prom_inst_0.INIT_RAM_0E = 256'h010C102229846300E969255860A82A20E0946489530362A1F57E0B271D34E114;
defparam prom_inst_0.INIT_RAM_0F = 256'h50B1E455099D4CACEC04830009954B427D34EF89444400004E65094415F1D34E;
defparam prom_inst_0.INIT_RAM_10 = 256'h4B3352333329503604B6A41042C435F373A433488DD8C408591542E353221B93;
defparam prom_inst_0.INIT_RAM_11 = 256'h4C10052E2DCCD2DBE9A70A22758F1505716E66F19720451260882BFAB52AFA58;
defparam prom_inst_0.INIT_RAM_12 = 256'hEEBA20643E4EA6EC8025D8E2D80886B0A6E14E000061604FFEFFEB1A4F8AA75A;
defparam prom_inst_0.INIT_RAM_13 = 256'h1B04FF37638B6A1AC29B8438000185813E0AD26000298511572AC7DC2689F284;
defparam prom_inst_0.INIT_RAM_14 = 256'h011405F72323229CE5E9AAB2499A582ED05037466F7CC5A9CF01FC0C05D4824A;
defparam prom_inst_0.INIT_RAM_15 = 256'hADC54422221044B4EBCD447BAC76669ECD580885965D10442208AD390544DB62;
defparam prom_inst_0.INIT_RAM_16 = 256'h844B4D8000028ADBF4B8A88444420827A6DAF3511EEF1D33A337F200001456DF;
defparam prom_inst_0.INIT_RAM_17 = 256'h99690C6A8853F6596498CFD964320E5C986009A324F94001456DFBDC54422221;
defparam prom_inst_0.INIT_RAM_18 = 256'hD9D1CEE8104B524CF9ED46D9DFCFFD35A41305A0E5F3939913DFCF343F78298C;
defparam prom_inst_0.INIT_RAM_19 = 256'h692926084010A94484408482C802204268A2FA31131B9A6B020893486DA4E520;
defparam prom_inst_0.INIT_RAM_1A = 256'h961426D2A68F4D924505B6C141046A3964B31693438DD3F0BB05F96BBEA804C5;
defparam prom_inst_0.INIT_RAM_1B = 256'h083FEFD2FDACF1A4218BF26FAD15604154121BFEF1FFC6739CF6D1A16B353024;
defparam prom_inst_0.INIT_RAM_1C = 256'h1E612C003AD38FAF06E2820B905186BA0D5528918658018516E92AB639150641;
defparam prom_inst_0.INIT_RAM_1D = 256'hE066494E69E524249A313A00DB4B163D172C000B1BCD76BB59316530101ABBB4;
defparam prom_inst_0.INIT_RAM_1E = 256'hD26ED2C8246059A64F365B236235D7A08AE61EA3319612816505A2281793445C;
defparam prom_inst_0.INIT_RAM_1F = 256'h8836722438EF4EC23B5B5A4CA991B9CC98098812012397FABF44468261BDF305;
defparam prom_inst_0.INIT_RAM_20 = 256'h6658D1B22763DC0E19176C7801EAC4B2C11582A2959800E4418D852B525200CC;
defparam prom_inst_0.INIT_RAM_21 = 256'h0B08C68809C843A084E8220E95630845A12B982CD9205980015268EC2BD3A015;
defparam prom_inst_0.INIT_RAM_22 = 256'hA29B55368A6D54DA29255248A55E19112E9BCC3DECD4938B7E2CA688C2815220;
defparam prom_inst_0.INIT_RAM_23 = 256'hD6907A96A494AB649149B24AAC9229255248A49549229B55368A6D564419258D;
defparam prom_inst_0.INIT_RAM_24 = 256'h9BDCA05430D247080E548C36D300C7C25E60C3C19874349434905E0AB5A004A0;
defparam prom_inst_0.INIT_RAM_25 = 256'hB6AB5625010811015FFA8051AF49D23F500CF708212C993925F07042592262E3;
defparam prom_inst_0.INIT_RAM_26 = 256'h00410000008242424937216602ACC05598312312896384884B1816603B2D3BF3;
defparam prom_inst_0.INIT_RAM_27 = 256'hCE610E93B7CB437EDAE9F2C951E20830000C50430C1041041040000000000000;
defparam prom_inst_0.INIT_RAM_28 = 256'h7FC6BE6DFF9AFB77FE6BECDFFCAFA9FF87FE59FFDFFFEBFFEFA208BAC4CE624D;
defparam prom_inst_0.INIT_RAM_29 = 256'hC8C33F840D95000000F4003FF0FFFDFFF0DFBFBABFB0BFA077F8A7FFFFF7FFD7;
defparam prom_inst_0.INIT_RAM_2A = 256'h5A03100A81523653B196AA2D3A4551A052D2C9A0D12882171931E030DD26999F;
defparam prom_inst_0.INIT_RAM_2B = 256'hAAAAAA0A00000000100000000000000000000003302A2088D342E8A3B6459107;
defparam prom_inst_0.INIT_RAM_2C = 256'h01123232323323333333333323234467545444444444567677667666AAAAAAAA;
defparam prom_inst_0.INIT_RAM_2D = 256'h3C001F803E441F8878983C700E0007000E000380033201010101010101010101;
defparam prom_inst_0.INIT_RAM_2E = 256'h0FC838001C000E0007000380038000E000E0003E600F9803E600F9803C001F80;
defparam prom_inst_0.INIT_RAM_2F = 256'hF67FFA9F7FCF9FD75FC553DEAAFFEAFD7FF7F7F7F7F7F7ADD7EB79883CE01E32;
defparam prom_inst_0.INIT_RAM_30 = 256'h8CCC8B55554CD8E7AFEBF5FAFD7EBF5F3E75EBF77AF8E1EBD79F3FAEBFED63DF;
defparam prom_inst_0.INIT_RAM_31 = 256'h00000000000000000000015FFEBAFD2EBFE974BBF7B5FFFFF6030FB55D4888CC;
defparam prom_inst_0.INIT_RAM_32 = 256'h80007FFF9C3F9C3FFFFF80007FFFFFE47FE57FFF91FFD1FF8000000000000000;
defparam prom_inst_0.INIT_RAM_33 = 256'h80002AAA800028782878114451FF80007FE411E47FFFD1E57FFFFE967E967FFF;
defparam prom_inst_0.INIT_RAM_34 = 256'h80002AAA9AAA9ABE1ABF9AAA9AAAAAAA80002AAA9EAAFEAAAAAE000007828782;
defparam prom_inst_0.INIT_RAM_35 = 256'h2AAE0000078811551145078800000000000002780278000011FFFFE451E43AAA;
defparam prom_inst_0.INIT_RAM_36 = 256'hAFFA80000000000000002AAA9ABFAAAA9D561D561D561AAA80001AAA9ABF9ABE;
defparam prom_inst_0.INIT_RAM_37 = 256'hECABEAABFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000007FAFFAFF;
defparam prom_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000007FFFFFFFD5552AAA;
defparam prom_inst_0.INIT_RAM_39 = 256'h1D5600001ABE2AAB800000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3A = 256'h1887000056180000280000007FFFFFFFFFFFFFFFFFFFFFFFEEAAABED8000AAAE;
defparam prom_inst_0.INIT_RAM_3B = 256'hA8002AAA80007FFF80000000019955AF819955AFE18001E3800000005AC60000;
defparam prom_inst_0.INIT_RAM_3C = 256'h0000788700000000088AEED56755555555555554D5062B587FFE801AB377AAAA;
defparam prom_inst_0.INIT_RAM_3D = 256'h07E6F8002FAF800007CA80000EBE000000008000000007E6000066BE000066BE;
defparam prom_inst_0.INIT_RAM_3E = 256'hFFF017FE5FFFF01FFF507FE3EFFF00001800012001D676BE01D680002FAF8000;
defparam prom_inst_0.INIT_RAM_3F = 256'hFF43FFF3F7FE3FFFF3FFFF3F7FE3DFFF41FFF7E7FE4AFFF40FFF7E7FE6AFFF3E;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[30:0],prom_inst_1_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 1;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hE3DFFF41FFF767FE4AFFF3EFFF017FE41FFF7EFFF727FE40FFF7EFFF6A7FE3EF;
defparam prom_inst_1.INIT_RAM_01 = 256'h000000000000000000000000000000000000000043FFF3F7FE3FFFF3FFFF3F7F;
defparam prom_inst_1.INIT_RAM_02 = 256'hAE2AAAFFFF800000007FFF81F800000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_03 = 256'h1F2CD72AAAAAAA9F807FFF806066607FE00000000000000000000000002AAAAA;
defparam prom_inst_1.INIT_RAM_04 = 256'hFAAAD5555555552AAAD535D554D506AAAAAB582AAAFFFE87FFAAAA801AACD700;
defparam prom_inst_1.INIT_RAM_05 = 256'h557FFF81085508000000002AAAD554AAAAAAAAAAAAAB5854AAFF52EED567557F;
defparam prom_inst_1.INIT_RAM_06 = 256'hFE2078000000007FFFFFFE00007FFFAAAAA8002AAA80007FFFDE405E557FFFD5;
defparam prom_inst_1.INIT_RAM_07 = 256'hF807D500007FFF800180001FFFCAAF80007FFFEAAA800000007FFE606600007F;
defparam prom_inst_1.INIT_RAM_08 = 256'h552AAA80007FFF80007555000000004AAA807A8000001E200620067FFE000075;
defparam prom_inst_1.INIT_RAM_09 = 256'h1F8000001F8000800000001FFFFFFF807AFFF87FFFA00660067FFE7FFE7FFFD5;
defparam prom_inst_1.INIT_RAM_0A = 256'hCF7FFFFFEAD7FC99FE7B77FFFFFFCDBFEE473FEA67FCF6FDC8CD95BF5FFFFF80;
defparam prom_inst_1.INIT_RAM_0B = 256'h040000AAB6DAAB2DAAEDA952AABFFFF000007FFFFEDB2AC9F61D9345FFFFFAC6;
defparam prom_inst_1.INIT_RAM_0C = 256'h4000040000FFFFFFD5AFC0701E3F8FFFFFFAAA002A2001A000041080C0080200;
defparam prom_inst_1.INIT_RAM_0D = 256'hCDAA402024ADAA4020A4160843FF040000400004FDFE4ADAA4020A40B0841FF0;
defparam prom_inst_1.INIT_RAM_0E = 256'hFF841BB840AA840EE84082840560407C040000400AD40000BFFFF400004FDFE4;
defparam prom_inst_1.INIT_RAM_0F = 256'hAC4F0F840000400AF40000BFFFF5FFFF40607406054060740009408D841FF041;
defparam prom_inst_1.INIT_RAM_10 = 256'hF5FFFF40607406054060740009408D841FF05FBFF5BB774A9554E9DD40905498;
defparam prom_inst_1.INIT_RAM_11 = 256'h0000023FC003FC0FFE0EFFFFFBFE1FDFF785FF7FB80FFBFEFFFFE01005FFBFFF;
defparam prom_inst_1.INIT_RAM_12 = 256'h4C00878008FC208DC3885438874388040884C0087800813208000080001FFFFF;
defparam prom_inst_1.INIT_RAM_13 = 256'hFFCFDFFCE5FFC81FFCFDFFCFDFFC7DFFC7FFFE8FC088DC388543887438804088;
defparam prom_inst_1.INIT_RAM_14 = 256'hC1B6DBF86FFE7FFFC7FFFC7FFFC7FFFC7BFFC83FFCFDFFC95FFC7DFFC03FFC83;
defparam prom_inst_1.INIT_RAM_15 = 256'h07FC0DB00FC00DB003F3FC007FBFFC3BFFC1B6DBF0000000000C007FBFFCDBFF;
defparam prom_inst_1.INIT_RAM_16 = 256'hA7F00555730C05557428403C70000000000000EAC03000EB000DCFFFFF5FFB00;
defparam prom_inst_1.INIT_RAM_17 = 256'h703C0ADDDF03FADDD03C0C3000FFF0000000000005FF5FAAA00000000FF5FFAA;
defparam prom_inst_1.INIT_RAM_18 = 256'hA000C03AA03ABF3AA000C000000000000EAB5000000D5AAD70F0000000355AAD;
defparam prom_inst_1.INIT_RAM_19 = 256'h00FC0D5FC03F000000000FC000000000003C700F03EACA950A550C000F000F3A;
defparam prom_inst_1.INIT_RAM_1A = 256'h1000000000AA0AAA00000A29600005570C3000D5C4440FFF80000000003FF020;
defparam prom_inst_1.INIT_RAM_1B = 256'h07C005C1C0000002A0030303F55FF5FD5EAB5EB005550AAAAE8000000AAAA200;
defparam prom_inst_1.INIT_RAM_1C = 256'h00000222200AA0000F3AA003C0003EAAB3C000000FEB7A57A140007F56010000;
defparam prom_inst_1.INIT_RAM_1D = 256'hF387F0EAB6AB0595755550000303FFC003EACEAABC0FC00005F5555C00000AF0;
defparam prom_inst_1.INIT_RAM_1E = 256'h0F00003C7000FDD55C00057DBFD2C0000387FFFFFFD2CFD2CFFFF387FFFFFFFF;
defparam prom_inst_1.INIT_RAM_1F = 256'h000003FC03CA0AA203C000000EFAC2AAAAD573FC03C253C165FF0D9550003C30;
defparam prom_inst_1.INIT_RAM_20 = 256'h0000000000000000000000000003700000370C015008280800F000000AAAA00F;
defparam prom_inst_1.INIT_RAM_21 = 256'h0000000000A0000000002FFF000000000000000000EAB6AB00000FF000001000;
defparam prom_inst_1.INIT_RAM_22 = 256'h2A0E08045008C4802EE80000000003D54200000A208080000220000000000004;
defparam prom_inst_1.INIT_RAM_23 = 256'h28C0282012C00A290292008880580AE08884400828C6EAA0824A10082848A2AA;
defparam prom_inst_1.INIT_RAM_24 = 256'hE64934B20B7FBBBBBBBBEAFA36AA360A00000000000000000000A8C820284862;
defparam prom_inst_1.INIT_RAM_25 = 256'h82DF4E5E006BEFAD82BEFA9294DB6DB77080006D27BF856F7BDFB6FFE924B2CF;
defparam prom_inst_1.INIT_RAM_26 = 256'h7035980857D4857D63BBFFCFFC94CC33EA0A08AFA67E5294AC777785F6FDA0AA;
defparam prom_inst_1.INIT_RAM_27 = 256'h05F11AFBCBCC4F8F8C55F79780000000000000720AE0C4D9B47AAFAB0AFA6777;
defparam prom_inst_1.INIT_RAM_28 = 256'h67BDEF3730C5041511430F1383A0C3C57A83DE250C502C054382800E5C5F863B;
defparam prom_inst_1.INIT_RAM_29 = 256'hBD34D2F2B0D0504AB6DB6DB841FC1CA9ECC80D103465550326F6F7BC9A5FB31D;
defparam prom_inst_1.INIT_RAM_2A = 256'h7777777777776555775C6AC5394EC4E061553DDDB1911792E9F6392BFD34D2F2;
defparam prom_inst_1.INIT_RAM_2B = 256'h99AD802E143AAEB8EA7957F137EFDE6A7924FA9B6DB6DB6DF7DF7DE0BB7C122B;
defparam prom_inst_1.INIT_RAM_2C = 256'h088801BC45494289BB3824A8EC1395EDB79806914912C97F3C3DFBF228A9FFFF;
defparam prom_inst_1.INIT_RAM_2D = 256'h39CE739CE548001E04771BCE5593A650054C49D3865554C90B374011702232A0;
defparam prom_inst_1.INIT_RAM_2E = 256'h01B5262AAA01FF5337081816840FFAEEBABBBEBFEFBFA500444EBFD50BA17E0B;
defparam prom_inst_1.INIT_RAM_2F = 256'h00FE1FE009FF1560AC008010022AE089012AA04255801BD60002100084004874;
defparam prom_inst_1.INIT_RAM_30 = 256'h0004102000012804A002010400000020000000640000000000000000024C40B5;
defparam prom_inst_1.INIT_RAM_31 = 256'h042448110820DA083002512108846891084219B6D42DFBA80020000002000000;
defparam prom_inst_1.INIT_RAM_32 = 256'hEAA8000FFFF36A8FFF0AA35200000001A82A420A000000000D04140129880021;
defparam prom_inst_1.INIT_RAM_33 = 256'h0440408808110004086000408100C0008102008102181020B020102181020BBC;
defparam prom_inst_1.INIT_RAM_34 = 256'h0081008100810204320A1028400810200400880811B401905081420040810020;
defparam prom_inst_1.INIT_RAM_35 = 256'h0006C0000000000000000953F7DF6444B000000254FDF7D80081008100810081;
defparam prom_inst_1.INIT_RAM_36 = 256'h5560301415580C00A832AB0180A055580C01807FCBDFDFFC49ED001800100014;
defparam prom_inst_1.INIT_RAM_37 = 256'h088442160E160E160E30650B070B070B071826F293C00060301E000301803506;
defparam prom_inst_1.INIT_RAM_38 = 256'h1084242108684214210822010010E2366648C42945614C2997B3333330884411;
defparam prom_inst_1.INIT_RAM_39 = 256'h288421084510842108821084211FFFE42108421090842108420410842108F67B;
defparam prom_inst_1.INIT_RAM_3A = 256'h080083F0B882102084368084105202002080F02120421A404004141040400410;
defparam prom_inst_1.INIT_RAM_3B = 256'h5554821084211ECF62190C43430402002199517FBDEF74042001087A02104148;
defparam prom_inst_1.INIT_RAM_3C = 256'hFCDB336CCDB33222226889A221A22226889A221911113444D110D50F7FF95555;
defparam prom_inst_1.INIT_RAM_3D = 256'h044444444444444000011110000044440000308888C56C56D86A53FDEF77F5DF;
defparam prom_inst_1.INIT_RAM_3E = 256'h19555422040804020BEF3AF3AFB38018F50E621CC21CD4060000000000000028;
defparam prom_inst_1.INIT_RAM_3F = 256'h003B00000000001121001121AA829080402000005555081210080433AAA80000;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[30:0],prom_inst_2_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 1;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'hFFFFFFFFFDAC4C91813646002C919106CCD1200503FFFFFBFFF1CDFFFFFFFD05;
defparam prom_inst_2.INIT_RAM_01 = 256'hB3A028195ADB49B49B49B49B40E2A3581D0F7FCD9B15E000028D83F0C880B8D2;
defparam prom_inst_2.INIT_RAM_02 = 256'h3CA692481FBF922AAC444E748F38B85C05B80AE17717F7092720C056A815D00A;
defparam prom_inst_2.INIT_RAM_03 = 256'h9236C3B20805C69AAA0206C40DB06CC5C4DB61DD7D5AC2F4E3BB05BF287981AF;
defparam prom_inst_2.INIT_RAM_04 = 256'h598C2C02A9DA923310C8C89236A48C99AC31ECA03111B393BC1B80C9AD264CEE;
defparam prom_inst_2.INIT_RAM_05 = 256'h930F4144695531DE12224A04D2604622208309401CC43310659C8393324C4294;
defparam prom_inst_2.INIT_RAM_06 = 256'hA0B16E48C06AE17041446E7B4806464931DE11E4C0C52EC08089252617611286;
defparam prom_inst_2.INIT_RAM_07 = 256'h000EC5455A4EE464734860B0C5325914C984D8620984D0C1625264E000088883;
defparam prom_inst_2.INIT_RAM_08 = 256'h8991B59444400000899C45800063332369B49A183029AED0882A0B08A1340000;
defparam prom_inst_2.INIT_RAM_09 = 256'h9A027FCF0C76330CA4899252492C1292264038BD030C8FF48308129261D684A4;
defparam prom_inst_2.INIT_RAM_0A = 256'h756D52CD2DA41A166C2133A0060EE72524CC129218C94913204A487D49491324;
defparam prom_inst_2.INIT_RAM_0B = 256'h84042A95D9957491AA000D7E804A628997212665934082016712BE083E2FB704;
defparam prom_inst_2.INIT_RAM_0C = 256'h861CB296049F0808247A822566B76A9C9364CEC384EC49A18C8D042155DD9C99;
defparam prom_inst_2.INIT_RAM_0D = 256'h379B90D3D99B925AC0DB024C125264699535476C34EE69A69199323795699749;
defparam prom_inst_2.INIT_RAM_0E = 256'hF89009C4C6525B3724B181B7849824A4C8D22A4A8ED869DC934C0332F5B12F88;
defparam prom_inst_2.INIT_RAM_0F = 256'h81A2476D4293624C2CB64CDB644D31102400234015115155113C44C24C2F5B12;
defparam prom_inst_2.INIT_RAM_10 = 256'hB56581C09C070C949A3537A98CC6A4C8482B018C6159204C91DB50A4D89A0424;
defparam prom_inst_2.INIT_RAM_11 = 256'h60DAB18B01604409A00153B3DEE458585A4B491050AC03120E449B27B9A501AF;
defparam prom_inst_2.INIT_RAM_12 = 256'h1321B705E5817411F5B377AEC1B1194B332A7B54D30697620820B06C66EDDC2C;
defparam prom_inst_2.INIT_RAM_13 = 256'hD827B40DDEBB0C652CCCA9ED534C3A5D9B916306558CA9D9DDFB7321B04F40D9;
defparam prom_inst_2.INIT_RAM_14 = 256'h61899A21CDB23216B734AA5F83A2A3352CFE09BD365051900380FC0FFB71B9DE;
defparam prom_inst_2.INIT_RAM_15 = 256'hD2523323231667DA048C26A4D299D30D85D39CBA5AAB98F73208E68BCE5A510C;
defparam prom_inst_2.INIT_RAM_16 = 256'hC479A30000006414DB4A46646462CA3ED1812319AD3426D4DC9B6000000320A4;
defparam prom_inst_2.INIT_RAM_17 = 256'h4F83DD82E9E0605005080181520144C94F972D15F9CA8000760A6D2527723239;
defparam prom_inst_2.INIT_RAM_18 = 256'h015A004047B010300026787810010730AB1A7CD69C042047A30E11321C20F2CD;
defparam prom_inst_2.INIT_RAM_19 = 256'h4C9594F9E35750613F4E523356E7A7290E72A52D11199E45D12EDA1D240002F4;
defparam prom_inst_2.INIT_RAM_1A = 256'h3ACFA4139A2C49B0098724AA5CEF4706D369BE96666860C66C8FB1ACDBA82C16;
defparam prom_inst_2.INIT_RAM_1B = 256'h35B29020920C028AF19D4042319784E19C8649D7E7DFED7E000274DB170C9011;
defparam prom_inst_2.INIT_RAM_1C = 256'h7BC1DAD6C8A85004EAFE0A4A523106228ED31AD7FDB5A8F62977A684313F95AA;
defparam prom_inst_2.INIT_RAM_1D = 256'h3F9BF3B9304992D647F68BCD68830F01CEDAD64780A0502010B009873972BB03;
defparam prom_inst_2.INIT_RAM_1E = 256'h4908508495AFA241700885BDF0E2581B4CDDC066FAC18C8CDC9C3B9B91893241;
defparam prom_inst_2.INIT_RAM_1F = 256'h7F5801C34B20808B8B2A2A20191800272198114A5A32694D2DC774AB0D012869;
defparam prom_inst_2.INIT_RAM_20 = 256'hD0FC59A31D82B530998C28C1492EC4338A162DF42CD842664D84973212FB2620;
defparam prom_inst_2.INIT_RAM_21 = 256'hCF6CC4CCA8506ABD1A05185C9CDBBD66A438003643DA91BB26A0C845C70F3E69;
defparam prom_inst_2.INIT_RAM_22 = 256'h46049C093812302460D9C1B382D2F0FABAC827C43E8CC20F29FDC664ACC071F9;
defparam prom_inst_2.INIT_RAM_23 = 256'h3819E484A126E2012705009188246049C09381230246049C09381232B46AA102;
defparam prom_inst_2.INIT_RAM_24 = 256'hB2B5EC5FBC5E661CE240F496E9580B888701DBF381C6232620D190E5852F36B2;
defparam prom_inst_2.INIT_RAM_25 = 256'h464FBEC6B661877D8088EA0891605E915D44AD5B94A4D4E97955D72909A64DA6;
defparam prom_inst_2.INIT_RAM_26 = 256'h10000000008242420DD11A9066520CCA41B6BF61C0F01245E47BE88F040CC260;
defparam prom_inst_2.INIT_RAM_27 = 256'h013AC2008323F01209A0C0F078C20030000C1045045041145040100104184106;
defparam prom_inst_2.INIT_RAM_28 = 256'h7FCBBED5FF9EFCD7FE3BF65FFCEFCD87F601E9CFCF83B3C7D68324B25A013BB0;
defparam prom_inst_2.INIT_RAM_29 = 256'hD8111FB04017000001FC0060FDFC7F703B20509E909E9FBFB7FD28007FF7FFC5;
defparam prom_inst_2.INIT_RAM_2A = 256'h78333126E1E67FE784FB02241B49C80CC1010879230DE61F9D13F27D8F64008F;
defparam prom_inst_2.INIT_RAM_2B = 256'h000000500050500010000000000000000000000A82AA4DAC9A24420BBE488417;
defparam prom_inst_2.INIT_RAM_2C = 256'h1013322322332222222222222332766777666776767674545445454455500000;
defparam prom_inst_2.INIT_RAM_2D = 256'hCBBBA7FFC9BBE4779767CB8FF2EE798BF2777CA3FC0100011001001100110011;
defparam prom_inst_2.INIT_RAM_2E = 256'hF237CFFFE7FFF3FFF9FFFCFFFCFFFF3FFF3FFFCFFFF3FFFCFFFF3FFFCBBBA7FF;
defparam prom_inst_2.INIT_RAM_2F = 256'h3BB13A877CC9E369A0E6414732627FC8291199119911F4D069349677CB1FE5CD;
defparam prom_inst_2.INIT_RAM_30 = 256'h40400799999100F8B120C04034100DA78E962C608B1A264C8193C6D3419DE146;
defparam prom_inst_2.INIT_RAM_31 = 256'h0000000000000000000001E71B4036800D00500B9AE1FF200BFDF45669840040;
defparam prom_inst_2.INIT_RAM_32 = 256'hFFFFFFFF9C3FF23FFFFFD5557FFFFFE47FE17FFF91FFC1FF8000000000000000;
defparam prom_inst_2.INIT_RAM_33 = 256'h80003AAA800038783878114451FFD5557FE411E47FFFC1E17FFFFE967E8DFFFF;
defparam prom_inst_2.INIT_RAM_34 = 256'h80002BAE9BAA9BBE1AAF9AAB9AABBABAFFFFBABA9EBAFAAEAAEE000007828782;
defparam prom_inst_2.INIT_RAM_35 = 256'h3ABE0000078811551141078A00000000000002780A78006011FFFFE441E42AAE;
defparam prom_inst_2.INIT_RAM_36 = 256'hA6BA020802880AA800002BAE9AAFBAAA9D561D561D561BAE80001BAA9AAF9BBE;
defparam prom_inst_2.INIT_RAM_37 = 256'hEAB3ECCBEB2B2B337551F555EAABF555E001EAABEAABACB3800A00026BA6BA6B;
defparam prom_inst_2.INIT_RAM_38 = 256'h0802002802A80288000A02800280028002880828000002A86CABFFFFD5552AAA;
defparam prom_inst_2.INIT_RAM_39 = 256'h1D5600001BBE3AAB82A80AAA082800AA08000000028002AA0AAA0A8802A80002;
defparam prom_inst_2.INIT_RAM_3A = 256'h1A07000017E4000028000000555575555555E001E00060006FAEF9F58000AAEE;
defparam prom_inst_2.INIT_RAM_3B = 256'hA8002AAA80000000080208027E18AA7FFE186E7FE1E019EBE780000056180000;
defparam prom_inst_2.INIT_RAM_3C = 256'h00007A1982A02AAA888AEEB5665555555555552AD418341F888B81EAB377AAAA;
defparam prom_inst_2.INIT_RAM_3D = 256'h7866F800567F80001FCA80000FFE07FF87FEE00000067866000066BE000061FE;
defparam prom_inst_2.INIT_RAM_3E = 256'h7FE817FEDFFFFBF7FEB07FEC0FFF84001FE0032001D655FE7F5760002E7F8000;
defparam prom_inst_2.INIT_RAM_3F = 256'hFFFD7FEBF7FEBFFFFBF7FEBF7FEC1FFF817FEFF7FEDDFFFBE7FEFF7FEDDFFFC0;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[30:0],prom_inst_3_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 1;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'hEC1FFF817FEEF7FEDDFFFC07FEFF7FE81FFFFF7FEE57FEBEFFFFF7FEDD7FEC0F;
defparam prom_inst_3.INIT_RAM_01 = 256'h01003F3A01211E121A3E1E1A031818181A26001E7D7FEBF7FEBFFFFBF7FEBF7F;
defparam prom_inst_3.INIT_RAM_02 = 256'hAE3ABAFFFFFFFF8001F55386AE2200002303213F0F1F0118262E061E3F3F2021;
defparam prom_inst_3.INIT_RAM_03 = 256'hF72CD72AAAAAAAFFE0606001807FE000607FFF87E01E601FE0000000003AEAAE;
defparam prom_inst_3.INIT_RAM_04 = 256'h57AAAB555555552AAAD54B552AD41AEAAAB41FAAAAAAAB87FFAAAA81EAACD701;
defparam prom_inst_3.INIT_RAM_05 = 256'h007FFF81080008000000004AAAD5552AD4D4AAAAAAB41FD4AFF6AAEEB5665555;
defparam prom_inst_3.INIT_RAM_06 = 256'h002018000000007FFFFFFFFFFF80002AAAA8002AAA80007FFFDE405E007FFF80;
defparam prom_inst_3.INIT_RAM_07 = 256'h5E60757FFF80006001800007AACAABFFFF80006AAA800000062006781E7FFE00;
defparam prom_inst_3.INIT_RAM_08 = 256'h552AAA80007FFF80007FFF800000007FFF81FF800000007FFE7FFE7FFF800075;
defparam prom_inst_3.INIT_RAM_09 = 256'h078000000780008000000007FFFFFF81FFFFE07FFFFFFE18067FFE7FF87FFFD5;
defparam prom_inst_3.INIT_RAM_0A = 256'h1CFFFFFFCCA7FDC9FE44E1FFFFFFC6FFE569BFBF27FC89FCAD5A938DEFFFFF80;
defparam prom_inst_3.INIT_RAM_0B = 256'h080000F3FFF736396CF1C6634C3FFFFFFFFFFFFFFAADD7F95EAC52EDFFFFF9EE;
defparam prom_inst_3.INIT_RAM_0C = 256'hC000080000FFFFFF994FFFFFFFC7F18000053C00F3210D3000C0101CF04CC400;
defparam prom_inst_3.INIT_RAM_0D = 256'hC7FECFFFCCFBFADC004C2AB8C4000C0000C0000DFDFCCFBFADE004C15E8C2000;
defparam prom_inst_3.INIT_RAM_0E = 256'hFF0C0BE8C1FF0C0FA8C3030C03A0C0800C0000C00D380000C000040000DFDFCC;
defparam prom_inst_3.INIT_RAM_0F = 256'h74D0100C0000C00D380000C00007FFFEC0607C0607C0605FE002C1808C2000C3;
defparam prom_inst_3.INIT_RAM_10 = 256'h07FFFEC0607C0607C0605FE002C1808C2000FF7FECB97DDF3FEDA9F5F0606C28;
defparam prom_inst_3.INIT_RAM_11 = 256'hFFFFF8C03FFC03F8000CFEEFE3FE1FDFF785FF78580FFDFEFFFFF01008004000;
defparam prom_inst_3.INIT_RAM_12 = 256'h1401880019F87985C718F8398D439980718140188001963798000100001FFFFF;
defparam prom_inst_3.INIT_RAM_13 = 256'hFFDFEFFDCAFFD7CFFDFEFFDFEFFD81FFF800009F8B185C718F8398D439980718;
defparam prom_inst_3.INIT_RAM_14 = 256'hBFF6DBFFAFFD7EFFD7EFFD7EFFD7EFFD82FFD02FFDFEFFDBAFFD80FFDFEFFD02;
defparam prom_inst_3.INIT_RAM_15 = 256'h0FD7CEB00DFFFEB00C3C0FFFBFB6DBDB6DBFF6DBFFFFFFFFFFFFFFBFB6D99B6D;
defparam prom_inst_3.INIT_RAM_16 = 256'hAF5F05DF300C05DF3C00433D70F0000F00000F6AC000C0EB0C0CCFFFF74D7B00;
defparam prom_inst_3.INIT_RAM_17 = 256'h7FC00ADDFCC03ADDFFC00C3C08FFF000C3FFC00004D74FAAA00000000D74DFAA;
defparam prom_inst_3.INIT_RAM_18 = 256'hA000303EA03FFFEEA0003000000003FFCBAB500000F5DAAD7F00000000F5DAAD;
defparam prom_inst_3.INIT_RAM_19 = 256'h13C005DC30D5C03FCC000DFFF00003FFC33D7030FFBACA950AA90C000FC0FFEA;
defparam prom_inst_3.INIT_RAM_1A = 256'h100150000AAA8AAA800038A9300005570C3C0035C44409D7A00000000007F121;
defparam prom_inst_3.INIT_RAM_1B = 256'h073C05C1C00022AAA000F0FC05DC05FD5FAB5EB0055509D7AA8000000FFFF211;
defparam prom_inst_3.INIT_RAM_1C = 256'hF00008080008A0000FEAA00C30003AAABC3000000FEB7A57A4700170DA300000;
defparam prom_inst_3.INIT_RAM_1D = 256'h7E47F0EAB6AB059FD555500000FC0DFFFFBAFAAAB3F00FFFF5F5555C00000FFF;
defparam prom_inst_3.INIT_RAM_1E = 256'h00FC033D700FDDF5D73C0F3EBFD2C0000387FFFFFFD2CFD1BFFFF387FFFFFD55;
defparam prom_inst_3.INIT_RAM_1F = 256'h05550CFF03C000021BC000000F0FCF0D08803CCCFFC25C3167F00D955000CC3C;
defparam prom_inst_3.INIT_RAM_20 = 256'h03FFC0C300FFC300C0FF00000003700000370FFFFFFFFFF3FF0000000FFFF33C;
defparam prom_inst_3.INIT_RAM_21 = 256'h000000000AA0000000028FFF23F3030000FF030F0FAAB6AB00000E40000013FF;
defparam prom_inst_3.INIT_RAM_22 = 256'h88082088822A0AA82A02000007F80F0008000008AAAAA000082000000FF00004;
defparam prom_inst_3.INIT_RAM_23 = 256'h0AA282AA2800A2A20AA0028280222800082020A88A08A028AA82AAA882A0A202;
defparam prom_inst_3.INIT_RAM_24 = 256'h0ADB64BEE783AFAFAFAFAAAA9D658EA50000000000000000000080A82088AA80;
defparam prom_inst_3.INIT_RAM_25 = 256'h9A35083C325A98D8BA29A65081AE9A6DF89111B1F282E89EF7BD6DA07B6DC100;
defparam prom_inst_3.INIT_RAM_26 = 256'h203FD4DFE97B2C5399017FCFFCAE58C4344EE68A732C62187B0202E34C3C5DB3;
defparam prom_inst_3.INIT_RAM_27 = 256'h93D236A7371494542AF14E2E200000000000000E060800197123DAF458A73020;
defparam prom_inst_3.INIT_RAM_28 = 256'hDF7BDEAC48189CD98D25E2F0F1507AA955F424B5081EDA76D83D4CB94E1D4F04;
defparam prom_inst_3.INIT_RAM_29 = 256'h801601E388C094DCFFFEDB609A35B073CA2350E1D29323A68D01EF7AF6FD44A0;
defparam prom_inst_3.INIT_RAM_2A = 256'h3222223633777003169B5305354DFFD0AD7361AF7F7F77CCD4C31DB8001601E3;
defparam prom_inst_3.INIT_RAM_2B = 256'h3A3A09CE9D0FCFC7FCE5B0053A74E9074FFC470D269349A49249248D9ED36EFF;
defparam prom_inst_3.INIT_RAM_2C = 256'h531C173F98D513B4C8B6D99050B63692FC3D2D4B8A3A55C061EE9D0239CA8044;
defparam prom_inst_3.INIT_RAM_2D = 256'h5AD6B5AD69080522CF7F948C6374F169B3DA7E278099998438CEADB7691B1BB0;
defparam prom_inst_3.INIT_RAM_2E = 256'h024F8C8CCCAB54C9A45DB240100EEEBEAFEBEEFFFBAABFEFBFF105015FFFC50B;
defparam prom_inst_3.INIT_RAM_2F = 256'h444302E54DFDBBF17E3CC118435540CDD7953194EFD75013108620010C10D8A0;
defparam prom_inst_3.INIT_RAM_30 = 256'hD55364A0A22F5AFD647BD13E82390EE8ADB165C064EB023135808A08A40C11F4;
defparam prom_inst_3.INIT_RAM_31 = 256'h3ABB6BE2BDC6913B993803F5FF95D1FDFD5F707DFFCE574100A2B15BBAAB1D55;
defparam prom_inst_3.INIT_RAM_32 = 256'hD555554AAAFF7EAEFF755CA8FAAFFAAA0D500D95C07F807FD0D646A407673D0D;
defparam prom_inst_3.INIT_RAM_33 = 256'hFB460C2942879C3A768002AE2A049AAF2831590E9DA0E9D907D8E9DA0E9D90FE;
defparam prom_inst_3.INIT_RAM_34 = 256'hC4385C38575E9D7B24F7E90A1DD5AB1F630C7D42870C212F9C1E7097A43EBFD7;
defparam prom_inst_3.INIT_RAM_35 = 256'h277117FD5575F57555755020E98E0EEE414A6CDC0818E9A8D77EDF7EDF7EC43E;
defparam prom_inst_3.INIT_RAM_36 = 256'hA8B85C2DEAAEB7580D08153E9F2FAA2954A92AFF637F7F7C795B75A5BF20412E;
defparam prom_inst_3.INIT_RAM_37 = 256'hD760099DB325B2050329009AC9B69196D996C01CE05FF5BD5EA3F82D6AB541B1;
defparam prom_inst_3.INIT_RAM_38 = 256'hC4210BD84287B0810EF6483AFCC404411005123FCF534B6D255DDDDDDD76B0AE;
defparam prom_inst_3.INIT_RAM_39 = 256'h2421084206EF7BDEF4D8C63B8C4D5553D84210840F7BDEF7BD70C631DC627BBD;
defparam prom_inst_3.INIT_RAM_3A = 256'hD7E625D1043087DC21408627EC8335F9895983085E10A066BF312C830EBF3122;
defparam prom_inst_3.INIT_RAM_3B = 256'hAAA8D8C63B8C4F77B82AF53D05D075F9883B79E3FEFF88210AD84282189FB20C;
defparam prom_inst_3.INIT_RAM_3C = 256'h1B6DDDB776DDDD88DCA332CCCA589D8B666D9992EC46D9994CCC9516D5550001;
defparam prom_inst_3.INIT_RAM_3D = 256'hF5DD775FF57DFDC9044F55524111D554AA6742ABFB3AB7AA002400E2F822E8A8;
defparam prom_inst_3.INIT_RAM_3E = 256'hA0020244810201E095D7F77DD7F6FFAF2472918404E42B33126EEC924C916D9C;
defparam prom_inst_3.INIT_RAM_3F = 256'h000B000000000007DEDDC7DE5548AF7FBFD99446AAAAB6A0AFF63B5F7FFED44C;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[30:0],prom_inst_4_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_4.READ_MODE = 1'b0;
defparam prom_inst_4.BIT_WIDTH = 1;
defparam prom_inst_4.RESET_MODE = "SYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'hFFFFFFFFFCA609110036440009911306CC853024F8FEFEFAFFF34DFFFFFFFA02;
defparam prom_inst_4.INIT_RAM_01 = 256'hE2DC354851FDB6492492DB6DB2C2B21BD10F5988910AC0000078BF43F88A03F0;
defparam prom_inst_4.INIT_RAM_02 = 256'hCC54D36B9B8794B8284CCE6F317D3A9C69B8D2EA770767196270810689A5D050;
defparam prom_inst_4.INIT_RAM_03 = 256'hDA2D55E2AA0EC7A6208246D41CB0E44E20B57302A8A7AA85D1442F9575FCFCF8;
defparam prom_inst_4.INIT_RAM_04 = 256'h11CC88A82890C22214C40052A43099B38C30DBB91919191316912289A5AECC62;
defparam prom_inst_4.INIT_RAM_05 = 256'h920694146A1F2494123083290B414632A28252205691A31867168311A04962D4;
defparam prom_inst_4.INIT_RAM_06 = 256'h00B5F70EE03F6A59141467F6AE48849324D491D4C0D5A88080C935A4A5457D06;
defparam prom_inst_4.INIT_RAM_07 = 256'h00266D571EE642023B8B6A3011321044C904D4634D06E2D47218410000088883;
defparam prom_inst_4.INIT_RAM_08 = 256'h8D25259666622224889F478952425B23E1F0EC1E2C354D3488A0812E05F08000;
defparam prom_inst_4.INIT_RAM_09 = 256'h8386800A492272EC308D249842A8B0C2349158DD4B4D3141C05D44C20D42AC30;
defparam prom_inst_4.INIT_RAM_0A = 256'h37FA1AA5BD244832E97E79F65352852184E9A0C250C8613A6A83095548613A41;
defparam prom_inst_4.INIT_RAM_0B = 256'h95065891911130B9A61211AE0398482992216225D8BADDBDF5529C3B144B250C;
defparam prom_inst_4.INIT_RAM_0C = 256'h964CB0C345218A4A298A2A0C443548BE916C44C184E449A10E8D86A55CCD1998;
defparam prom_inst_4.INIT_RAM_0D = 256'h331311D8DFD31678C8D5E2495353406B917446A8B4F44127B599726685B99248;
defparam prom_inst_4.INIT_RAM_0E = 256'h7EDBC8C4EC465FA62CF591ABC492A6A680D622C88D5169E8826E4B32C5B1A7EB;
defparam prom_inst_4.INIT_RAM_0F = 256'h83A14629CA022ACCCDFBF8FFBC09717C3F188B50404444404046C4961DAC5B1A;
defparam prom_inst_4.INIT_RAM_10 = 256'h7FDC0AC023AC1C04B827921B1C9424CA0A751144E910A0E8509A72048ABA1422;
defparam prom_inst_4.INIT_RAM_11 = 256'h60DAA19F9BF35D4BB8C51391AF447CECFCDF989050A4025B0E6C3AB7B5A5F3FF;
defparam prom_inst_4.INIT_RAM_12 = 256'hEDC3B24C4785A449A5B2B62CC3139D89B0A635579A0713638E38F82367EF7023;
defparam prom_inst_4.INIT_RAM_13 = 256'h58226F2AD8B3067626C298D57E681C4D9F911B06550C89C89A83A211B0C4F2DF;
defparam prom_inst_4.INIT_RAM_14 = 256'hCD9C9AFF4F1111084338AA0423F2231F59E271DC2DDCC195057E000002B5B0C6;
defparam prom_inst_4.INIT_RAM_15 = 256'hF87376011184219C0DEC227DF81D82BB8DD11C8A823F99E7118067098E1A1B4E;
defparam prom_inst_4.INIT_RAM_16 = 256'h421DC1000000CC95FE0E6EC02220C70CE0837B089F7C8780EC16E200000664AF;
defparam prom_inst_4.INIT_RAM_17 = 256'h108DA98ED1A2834434018A0D186A44DD11C52D0441E8C000224AFF0773201110;
defparam prom_inst_4.INIT_RAM_18 = 256'h2152820F99F4903490A95D210481FBA2A3500936BD25001883D097A221589860;
defparam prom_inst_4.INIT_RAM_19 = 256'h459980112BD16875966C441B45C336220472F60888008E4789ACD21C0C4295D4;
defparam prom_inst_4.INIT_RAM_1A = 256'h2B99341122036DF11D86B6C351474F07C3E1BADE67B078A6E88F314DBF820482;
defparam prom_inst_4.INIT_RAM_1B = 256'h2525AEB76DE9D78A79BE416E3583E0F1DC9703FDA37E966B504557AE00FC2541;
defparam prom_inst_4.INIT_RAM_1C = 256'h7F31F4078B36D037E8E602CA562524520C8212D599E80D0279660496A18795C2;
defparam prom_inst_4.INIT_RAM_1D = 256'h418BD3DC2B4196961B2433082AC65510DDF4066A8E8743A1D0A301823878A207;
defparam prom_inst_4.INIT_RAM_1E = 256'h09001401A52250615A4E025320B79E33EACA9246EBB684DCA98E19B8C581A711;
defparam prom_inst_4.INIT_RAM_1F = 256'h9D414A610188C78B0A2A2A293118A088A390399E58B3E87D0FD3669B05140028;
defparam prom_inst_4.INIT_RAM_20 = 256'h2AC859321B036D20108A68E94BA69432CA540E1065D2FCF309083B1B5BC7B42A;
defparam prom_inst_4.INIT_RAM_21 = 256'hE94AA0C42844F8950A05585C1C9BAC66A51A090951AA018904B0CED446CE3045;
defparam prom_inst_4.INIT_RAM_22 = 256'h047018E031C06380C7008E0114C04D3820E88864E408D3094B65846EA6ED4A73;
defparam prom_inst_4.INIT_RAM_23 = 256'hB818E4863C04455C0206EE01178047018E031C06380C7008E011C0226628A1B8;
defparam prom_inst_4.INIT_RAM_24 = 256'h9B6C7E8BAE8E0214C087943EE3104F4987F09B63BBC621862298984D11A37631;
defparam prom_inst_4.INIT_RAM_25 = 256'h7C8E5FB79440D94882728608104E1ECE50C4DB3B1102C0D921B3B62245864160;
defparam prom_inst_4.INIT_RAM_26 = 256'h000002082186424201851A2266444CC889B27A6A455436A96458940927182082;
defparam prom_inst_4.INIT_RAM_27 = 256'h04474380F2A00013C0B8A0001C441831041C51430C5141141140004100104100;
defparam prom_inst_4.INIT_RAM_28 = 256'h7FC3BF3DFF8EFE37FE3BFADFFDEFEB87E601DBCFDF83CFC7E68306A208054B55;
defparam prom_inst_4.INIT_RAM_29 = 256'h929115204017000001DC0060F0FC7CF03D807FF6FFFCFFC037FCF2007FF7FFE3;
defparam prom_inst_4.INIT_RAM_2A = 256'h583829AEF4A012A7411B8A2C1B4DDAACC1818DB1230CC61D1503F87F10F65A8A;
defparam prom_inst_4.INIT_RAM_2B = 256'hEEEEEB4EEE4E4EEEDEEEEEEEEEEEEEEEEEEEEEE0B423000EDB44480A22089014;
defparam prom_inst_4.INIT_RAM_2C = 256'h00032222222332323232323223336776666667776677676767766666404EEEEE;
defparam prom_inst_4.INIT_RAM_2D = 256'hCBBBA63FC9BBE4779767CB8FF3FFF9FFF3FFFCFFFC1100011110111111110000;
defparam prom_inst_4.INIT_RAM_2E = 256'hF3FFCFFFE7FFF3FFF9FFFCB37C9CFF2CDF273FC99FF267FC99FF267FCBBBA63F;
defparam prom_inst_4.INIT_RAM_2F = 256'hFFFF3567FCE1029148E023C7FFFE4048291199991111F4CE66331FFFCFFFE7FF;
defparam prom_inst_4.INIT_RAM_30 = 256'h000447E1FFFF8840D978E6523F9FCA454D193077CB93324C99C2052291EC03C7;
defparam prom_inst_4.INIT_RAM_31 = 256'h000000000000000000000147149229248F49748D9FDEFF2006030C379E444404;
defparam prom_inst_4.INIT_RAM_32 = 256'hD5557FFF9C3FC83FFFFF80007FFFFFE47FF87FFF91FF87FF8000000000000000;
defparam prom_inst_4.INIT_RAM_33 = 256'h7FFF80007FF828780078114451FF80007FE411E47FFF87F87FFFFE967E837FFF;
defparam prom_inst_4.INIT_RAM_34 = 256'h80002AAA9AAA9ABE1AAB9BAA9AAAAAABFFFFAAAA9EABEAAABAAE07FF87838780;
defparam prom_inst_4.INIT_RAM_35 = 256'h2AAE007F8788115511500782FFFFAAAAFF8002782878000011FFFFE407E42AAA;
defparam prom_inst_4.INIT_RAM_36 = 256'hFEBF8A0A0AAA0AAA00A02AAA9AABAAAA9D561D561D561AAA80001AAA9AAB9ABE;
defparam prom_inst_4.INIT_RAM_37 = 256'hF32BEAADEAB2B2AAF2A9F7FDEFE3F555E7F9EAABEFFBAAAB802A00026BFEBFEB;
defparam prom_inst_4.INIT_RAM_38 = 256'h082200AA0AAA0AAA002A0AA20AA20AAA0AAA08AA08000AAA6ACBFFFFD5552AAA;
defparam prom_inst_4.INIT_RAM_39 = 256'h1D5600001ABE2AAB8AAA0AAA08AA02AA080008020AA20AAA0AAA0A8A0AAA0082;
defparam prom_inst_4.INIT_RAM_3A = 256'h78998000667428002AAA80005555755555558001E00000006BFA81F58000AAAE;
defparam prom_inst_4.INIT_RAM_3B = 256'h280000AA80007FFF820A0A0A781954607818666039FF81EBF87E000017E00000;
defparam prom_inst_4.INIT_RAM_3C = 256'h1F8018E00AA80000088AEEAB7E555555555552AAD0605060088AFEAAB377AAAA;
defparam prom_inst_4.INIT_RAM_3D = 256'hF866B800666000019FFFF8007F801EBF9EBEFE800001F866000061FE00180180;
defparam prom_inst_4.INIT_RAM_3E = 256'hFFF7EFFF5F7FE3FFFF67FFF007FE6C001E1F9B0001D7D5807D577E8058600001;
defparam prom_inst_4.INIT_RAM_3F = 256'hFE7EFFF7CFFF7C7FE7CFFF7CFFF007FE7EFFF7FFFF7B7FE00FFF7FFFF7F7FE00;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[30:0],prom_inst_5_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_5.READ_MODE = 1'b0;
defparam prom_inst_5.BIT_WIDTH = 1;
defparam prom_inst_5.RESET_MODE = "SYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'hF007FE7EFFF77FFF7B7FE00FFF7EFFF7E7FE7FFFF61FFF007FE7FFFF7FFFF007;
defparam prom_inst_5.INIT_RAM_01 = 256'h1F213F3B09253F333F3F3F3F073D3D3F3F2F203F7EFFF7CFFF7C7FE7CFFF7CFF;
defparam prom_inst_5.INIT_RAM_02 = 256'hAE2AAAFFFFFFFF800075539AAE140C002707133F1F3F013D2F110F3F3F3F2033;
defparam prom_inst_5.INIT_RAM_03 = 256'hD72CD72AAAAAAAE06060607FE01F8001807FFF98187FF87FF8600000002AAAAA;
defparam prom_inst_5.INIT_RAM_04 = 256'hB52AAAD55555557AAAAD54D2AAD06ADAAAD06AAAAAAAAA87FFAAAAFEAAACD77E;
defparam prom_inst_5.INIT_RAM_05 = 256'hAAFFFF81082AA000000000552CD55553555554AAAAD06ACAFD7EAAEEAB7E554A;
defparam prom_inst_5.INIT_RAM_06 = 256'h00201E0000000067FFFFFFFFFF80002AAA280000AA80007FFFDE405EAAFFFFAA;
defparam prom_inst_5.INIT_RAM_07 = 256'h57F81F7FFF800078018000006ACAAAFFFF80006AAA8000000620063F807FFE00;
defparam prom_inst_5.INIT_RAM_08 = 256'h552AAAFFFF80007FFF800001FFFFFF800000007FFE7FFE000000007FFF800075;
defparam prom_inst_5.INIT_RAM_09 = 256'h000000000000009878000001D5755500004B804AAA8000060620067FE07FFFD5;
defparam prom_inst_5.INIT_RAM_0A = 256'h877FFFFFCF83FF1BFE1FA0FFFFFFEFBFEFF6FFEC6FFC3F7DFEE7C78777FFFF80;
defparam prom_inst_5.INIT_RAM_0B = 256'hF80000E3E39FC639EF3EFC7800C00007FFFFFFFFFEC15A60767F7741FFFFFFBB;
defparam prom_inst_5.INIT_RAM_0C = 256'h3FFFF00000FFFFFF9F07C0701D27498000063FFFCCDEFD3FFFFFEFEF0FB3FFFF;
defparam prom_inst_5.INIT_RAM_0D = 256'hFD3930001339392C00F3E777380073FFFF3FFFF3FFFF339392E00F3F3C73C007;
defparam prom_inst_5.INIT_RAM_0E = 256'h55F3EBF73E0073FAA73D2BF3FFDF3F01F3FFFF3FFCD00000FFFFFBFFFF3FFFF3;
defparam prom_inst_5.INIT_RAM_0F = 256'hFB206033FFFF3FFCD00000FFFFFBFFFB2060420604206041E00B3F3973C0073F;
defparam prom_inst_5.INIT_RAM_10 = 256'hFBFFFB2060420604206041E00B3F3973C00735EAB3E57E204002A7541AA57307;
defparam prom_inst_5.INIT_RAM_11 = 256'h0000003FC000000FFFFCBEFFFFFFFFDFF7FDE17FFFF7F9FEFFFFFFEFF3FFFFFF;
defparam prom_inst_5.INIT_RAM_12 = 256'h83FE703FE7AF0E7F3FE703F6753F66D7BE783FE703FE63F0E7FFFE00001FFFFF;
defparam prom_inst_5.INIT_RAM_13 = 256'hFFDFFFFDC3FFD01FFDFFFFDFFFFD00FFDFFFFF7AF1E7F3FE703F6753F66D7BE7;
defparam prom_inst_5.INIT_RAM_14 = 256'hBFFFFFFFDFFDF9FFDF9FFDF9FFDF9FFD01FFDFDFFDFFFFDF7FFD01FFDFDFFDFD;
defparam prom_inst_5.INIT_RAM_15 = 256'h07FEBEB00D7AAEB0000008923FBFFBBBFFBFFFFFFFFFFFFFFFF8923FBFFB7BFF;
defparam prom_inst_5.INIT_RAM_16 = 256'hA7FACF503C300F5033FFF03D73FCC03FC00005EACCF00FAB03030FFFF7FD7B00;
defparam prom_inst_5.INIT_RAM_17 = 256'hF0000FFD7FC00FFD70000F3FF8FFF000C3FFC0000FD7FFAAA3CC00000D7FDFAA;
defparam prom_inst_5.INIT_RAM_18 = 256'hA000003AA03FFFAAA00000000300C3FFCAAFF0000F55FAABF00000000F55FAAB;
defparam prom_inst_5.INIT_RAM_19 = 256'h0FAAA5FFD355C0FFC73C0D7AA00003FFC03D7F305FAAF9550A950C000FCFAFAA;
defparam prom_inst_5.INIT_RAM_1A = 256'h1AAA40000956A556A000DFFFC00005570F3FF00F04440957A000000005555020;
defparam prom_inst_5.INIT_RAM_1B = 256'h0C070705C00AAAA95000000005FFFFFD5EAFFFFF05550957AA8000000FFFD200;
defparam prom_inst_5.INIT_RAM_1C = 256'h50000222200A2002AFAAAF0C1000DAAAA03000000FEB7A57A00C05C0389C5000;
defparam prom_inst_5.INIT_RAM_1D = 256'h7907F0EAAEAB0FF50FFFF00000000D7AAFAADAAAA0000AAAAFF5555C00000555;
defparam prom_inst_5.INIT_RAM_1E = 256'hFFD7003D70F57D7F5FEB003EBFD2FFFFFF87FFFFFFD2CFD06FFFF387FFFFFDFC;
defparam prom_inst_5.INIT_RAM_1F = 256'hF000ACC3C7D5500200C000000EFADEF909803F3FFFFFFFFFFC0003FFF03FF33F;
defparam prom_inst_5.INIT_RAM_20 = 256'hC3FFC3C3C3FFC30CC3FFC00000FF70000FF70C3105C000000000000005555000;
defparam prom_inst_5.INIT_RAM_21 = 256'h000000000000000000080FFF23F3C30003FFC33FCFAAAEAB00000E40000013FF;
defparam prom_inst_5.INIT_RAM_22 = 256'hA28A8A8A20A2AA888220000002AFFD554000000A2000000002200000055FF004;
defparam prom_inst_5.INIT_RAM_23 = 256'hA088AA8028A0AAAA2A2200A02A2000AAA0200A2222AA828220A8A0A2008208A8;
defparam prom_inst_5.INIT_RAM_24 = 256'h76493638677BEEBBEEBBFFFFBBFEEFBE30993B350C4800000000A88A02A88AAA;
defparam prom_inst_5.INIT_RAM_25 = 256'hBF2D882D224A56541F254E52918E3864459919F5B69CC996B5AD24B06924BE5B;
defparam prom_inst_5.INIT_RAM_26 = 256'h50018123ED9A3E4ADBBAC000022A18964EE447C953786318515775D2CB4C59B1;
defparam prom_inst_5.INIT_RAM_27 = 256'h82C2329595109416B9F92A2B2000000001FFFFFFFFE8C889517BDB347C959577;
defparam prom_inst_5.INIT_RAM_28 = 256'hCB5AD625734C94D8CB85A320D5996ACA59D0E6B10C129810CB8CCF3DEF298F9C;
defparam prom_inst_5.INIT_RAM_29 = 256'h8395196A808490C6F6DA4920A3394A53B90CDDBBE6D6665B54C56B58DB6D3425;
defparam prom_inst_5.INIT_RAM_2A = 256'h333333332133311386194340B02CC54ECB33358DB1191054C32F99A86395196A;
defparam prom_inst_5.INIT_RAM_2B = 256'hAFBBCDCA0C8A82A02B88B3EAECD9B2086DB4E643A1D0E87471C71C719B58813B;
defparam prom_inst_5.INIT_RAM_2C = 256'h5B9BE5AC88CD9146D8C31197FF70B32A94BC28E2F1D645C3640B36FDB93F7F3E;
defparam prom_inst_5.INIT_RAM_2D = 256'h18C6318C610804D28F580F2C233FE838B2C87FA72ABBBA02692BCE484DD2F6AF;
defparam prom_inst_5.INIT_RAM_2E = 256'h842D8870F067983838D9DC00000FAFBAEEEFBEAAABEEFFFBAAEFEABEF045015B;
defparam prom_inst_5.INIT_RAM_2F = 256'h54BF15455C239470A604C01BBB75E08C23847174AADDDABB315C48069C21B944;
defparam prom_inst_5.INIT_RAM_30 = 256'h28A1AA579DB89B4931249A43B562F0C5CE37FF8D1A03E5EBC1F7F7FF78CD44B1;
defparam prom_inst_5.INIT_RAM_31 = 256'h815084084A8808C242A44C4040CA862142840331D41D03415B5003F04403E28A;
defparam prom_inst_5.INIT_RAM_32 = 256'hFFFFFFE55517950C54754CA105500552928000759F807F8014A8A14A20104241;
defparam prom_inst_5.INIT_RAM_33 = 256'hDA8810118302100000A4C08832405008304000800028000096D0000280000931;
defparam prom_inst_5.INIT_RAM_34 = 256'h9830183018200080469568801B902697D21A45830218003C885221D81B76F6DE;
defparam prom_inst_5.INIT_RAM_35 = 256'h312D55D7D777C8A228A221037FDFC000537D878040DF7FDFDB7680001B768036;
defparam prom_inst_5.INIT_RAM_36 = 256'hA81D0E886286A351848150D46A412201E0F08055E3F5F5D6D958202B5413141B;
defparam prom_inst_5.INIT_RAM_37 = 256'h176000D0D2A0D2A8D0020C2C695431D4300346284015FA1D0E81D7F868345090;
defparam prom_inst_5.INIT_RAM_38 = 256'h885AD216B4A00D6AD000254037285555444510E52E4528E1304CCCCCC960B000;
defparam prom_inst_5.INIT_RAM_39 = 256'h535A000008000000012028005000000006B400000B4000000022294002800301;
defparam prom_inst_5.INIT_RAM_3A = 256'h01B942A0134D6ACB5A537943284CC06E50A8ACD695AD29980DCA104C900DCA11;
defparam prom_inst_5.INIT_RAM_3B = 256'h0001202800500060314CA601B90A806E50C408A8000023DAD7FEB4ADE50CA133;
defparam prom_inst_5.INIT_RAM_3C = 256'h5F24CC93324CC8999896660CCA8CCC882220888864CCC33304446E300002A802;
defparam prom_inst_5.INIT_RAM_3D = 256'h0C6646664CCEE6595DC99336577064CDDC0054C8CB329328490043777FDD7F57;
defparam prom_inst_5.INIT_RAM_3E = 256'h282A882452B4BA5D0FD7D5FFF7547FA72072B9E44CE47F303659A4763FCCA402;
defparam prom_inst_5.INIT_RAM_3F = 256'h001400000000000800000AD6001C42140A004FFCAA22114869757A4455543B33;

pROM prom_inst_6 (
    .DO({prom_inst_6_dout_w[30:0],prom_inst_6_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_6.READ_MODE = 1'b0;
defparam prom_inst_6.BIT_WIDTH = 1;
defparam prom_inst_6.RESET_MODE = "SYNC";
defparam prom_inst_6.INIT_RAM_00 = 256'hFFFFFFFFFFA68F9782365E084CBDB9237451742582FAFAFAFFF864FFFFFFFA02;
defparam prom_inst_6.INIT_RAM_01 = 256'hA3BC2F0D9FB5B6DB6492DB6CB242B72823094C6C082AA000010BFF3F7BAA0B30;
defparam prom_inst_6.INIT_RAM_02 = 256'h5C071681291F15D2AC44C6E9974C1A0D60BAC0E83714664C232080068D81D810;
defparam prom_inst_6.INIT_RAM_03 = 256'h481BD1D1E72EE1242AAB620089844C66406E1A882000280DF957524AA87522D2;
defparam prom_inst_6.INIT_RAM_04 = 256'h550A1C4009AB426F3FB98C81B2D08F3D21B8B71D311991319499A098C404C47B;
defparam prom_inst_6.INIT_RAM_05 = 256'h0F4E8014625774FC9146DB6D4B2F0747B282DB68CE5D57A22E449111F04F8F72;
defparam prom_inst_6.INIT_RAM_06 = 256'hAA279502002508E1001467ED876282DB74FCD8BCC6D6A4C89C6976BE26264907;
defparam prom_inst_6.INIT_RAM_07 = 256'h00137A9F55525C4C788B6A137913BBE44B8E0E656B9E22D43A29EC20426AE8D1;
defparam prom_inst_6.INIT_RAM_08 = 256'h9DFE75B64752031C9889024A34E3C9308050FCCE1924CD2488AAA3B304409554;
defparam prom_inst_6.INIT_RAM_09 = 256'h91A6998E3D2277C4D08DFE684FA0134277F71FE8461896E4E26C73427DA604D0;
defparam prom_inst_6.INIT_RAM_0A = 256'h649254E5A0265AE162FFA0D144C4C826846F83425019A11BCE0D096C19A11BFA;
defparam prom_inst_6.INIT_RAM_0B = 256'h940AF895D7BFB7CB3E43454F07D8E02897222664A3B2DBFC9153999626000006;
defparam prom_inst_6.INIT_RAM_0C = 256'h924C84835086022084B32E4648CE8C1B9444CD45C45CD9838E82B9B2BC8DA6EB;
defparam prom_inst_6.INIT_RAM_0D = 256'hE3BD04889B5314D018E5FA3DD3D3E3813D27C4A0519427972082666785A287C9;
defparam prom_inst_6.INIT_RAM_0E = 256'hA64C2CCD54031EEE29A431CBF47BA7A7C7037A6F8940A3284F2F6104C184EA74;
defparam prom_inst_6.INIT_RAM_0F = 256'hC353863D5A475070456D24B69A1C4841090AE58064246642490E05CB684C184E;
defparam prom_inst_6.INIT_RAM_10 = 256'h7FE418508477AFB61EB453C9AC529693015002C58A69B0F4E09F5615D41D3946;
defparam prom_inst_6.INIT_RAM_11 = 256'h89988024188B10478857D1332940A626208450D7D6A787554456D2BCAC2561FF;
defparam prom_inst_6.INIT_RAM_12 = 256'hABD3336D4E43F2209084A606139B990385FA2513080E070FDF7DEC368DCC4076;
defparam prom_inst_6.INIT_RAM_13 = 256'hC2226BB2981844640C17E8946820381C3711B4444401E9999290A0198444BA1F;
defparam prom_inst_6.INIT_RAM_14 = 256'hDFBE7C962DE363308F080084D142B3125BA230541B8EC198408103FBF4A13074;
defparam prom_inst_6.INIT_RAM_15 = 256'h603E83F2633E6F84464023C9600541F7ABB154ACA2A4AF3BF389E11F987920DD;
defparam prom_inst_6.INIT_RAM_16 = 256'h66F8452AAAA917E96C07D07E4C678B7C22919008F6580300280DCA000008BF49;
defparam prom_inst_6.INIT_RAM_17 = 256'hCA4564C6B89A1E91E803E87A40F80659422620204C8A80008BF4B603A83F2633;
defparam prom_inst_6.INIT_RAM_18 = 256'h4D62425FCA192B260808AA1C404041963A5B5C8563108A4A0CBE4193A031406D;
defparam prom_inst_6.INIT_RAM_19 = 256'h393E36B18D95FF6D3882D673D5EC416B45509FFB9BB9160FB9841949DC94D094;
defparam prom_inst_6.INIT_RAM_1A = 256'h92ABC691F27E82484884924A9F15552100A041094BF3387468EB20C9B7AA8ED0;
defparam prom_inst_6.INIT_RAM_1B = 256'hB5D9ACB6C965E761E93A100073974207B8E474D4A15A84629401225320039335;
defparam prom_inst_6.INIT_RAM_1C = 256'h35352497F37E75BEDAF6034B5375EAF20EB339A7DE4928301B77E680701F0E4B;
defparam prom_inst_6.INIT_RAM_1D = 256'h068882701D5022508A931AC400404409CD2494620B0582C160C5D022A920F126;
defparam prom_inst_6.INIT_RAM_1E = 256'h0510250298EBE0206C04036CB06DE71546738954E16104293F4F139F1280E205;
defparam prom_inst_6.INIT_RAM_1F = 256'h2D12688181404045103830211009A8215113114A6813B2774BB678E8462D41A2;
defparam prom_inst_6.INIT_RAM_20 = 256'h6E2C29C192044A2282D3544D050602818863A275C2C5FF4086081B0C030ED04E;
defparam prom_inst_6.INIT_RAM_21 = 256'h6C166006EADD225028344D43CF60A2A64198810917D901E9969075ED46CF32C9;
defparam prom_inst_6.INIT_RAM_22 = 256'h8CB9097212E425C84B90972131444C5C9278218C320819E401B4744ECD6C2AF3;
defparam prom_inst_6.INIT_RAM_23 = 256'hBA68EC402E424BCE4245E7212DC84B9197232E465C8CB9197232E466A87E901C;
defparam prom_inst_6.INIT_RAM_24 = 256'hBC4D5529C5254C16C4936B4B3F7E2EE5266E48D09DE2068204A1CC47223A3253;
defparam prom_inst_6.INIT_RAM_25 = 256'h2019D1AA5304CA2C0143480D93465C6829031355B59E7C9162352B6B6CA60040;
defparam prom_inst_6.INIT_RAM_26 = 256'h103080080144424373F219E2667C4CCF89B3693804651264C53AF8258200E808;
defparam prom_inst_6.INIT_RAM_27 = 256'h414A248130C61094C088399CD8C20050001430C20861840450431071030001C4;
defparam prom_inst_6.INIT_RAM_28 = 256'h7FC2BF7DFF8AFD77FE2BF7DFFCAFC3FFD7FF97FFFFFFFFFFE78224928B400FAC;
defparam prom_inst_6.INIT_RAM_29 = 256'hE2491F84489500000134007FC5FFFDFFFF7F9F9F9F9A9F8037FDF3FFFFF7FFFF;
defparam prom_inst_6.INIT_RAM_2A = 256'h62F4E1ADE4244B32943032ED102E93B8A16149B5B20AC45296242088CF20938F;
defparam prom_inst_6.INIT_RAM_2B = 256'hFAFAFE5AFA0F5AFACFAFAFAFAFAFAFAFAFAFAFACB488201D190E0783A91C0F03;
defparam prom_inst_6.INIT_RAM_2C = 256'hCD03ABEFEF23AB2233223322BBAB7777777776666677777777777777005AFAFA;
defparam prom_inst_6.INIT_RAM_2D = 256'hDFFFAFFFD9BBEC77B767DB8FF6EE7B8BF6777DA3FDD0CDCCDCDCDCDCDCDCCDCD;
defparam prom_inst_6.INIT_RAM_2E = 256'hF637DB9DEC9FF6E77B27FDB37D9CFF6CDF673FD99FF667FD99FF667FDFFFAFFF;
defparam prom_inst_6.INIT_RAM_2F = 256'hFFFF7FEFFDEBF693FDC7DEAE006AC0582BBB33333333FDEAF57AB677DB1FEDCD;
defparam prom_inst_6.INIT_RAM_30 = 256'h404273E0000600FDFB79E6D27FB49A4D1C3F7EDD5C3362CD9BD7ED27FBED9EAF;
defparam prom_inst_6.INIT_RAM_31 = 256'h0E51B1B1B11111BB11BB114F3FFF7FAFDA497499B514FF6006030C3818677004;
defparam prom_inst_6.INIT_RAM_32 = 256'h80002BFF9C3F80FFFFFFFFFFFFFFFFE47FFFFFFF91FFFFFF90E91BB11BB11BB1;
defparam prom_inst_6.INIT_RAM_33 = 256'h7FFF80007FF828780078114451FFD1FFFFE411E47FFFFFFFFFEAFE967FA02AAA;
defparam prom_inst_6.INIT_RAM_34 = 256'h80007AAAFAAE9ABE7AAA9AAA9BAAAEAAAAAAAAAA9EAAABAAAAAE07FF87828780;
defparam prom_inst_6.INIT_RAM_35 = 256'h2AAF81FF87881155115507E07FFF80007FE0027801F8006011FFFFE47FE47FFF;
defparam prom_inst_6.INIT_RAM_36 = 256'hAE9A880208220AAA00A07AAA9AAAFFFFFD579D561D567AAAFFFF9AAE9AAAFABE;
defparam prom_inst_6.INIT_RAM_37 = 256'hEAADF2CBECAAAAB2F2A9F61DEEA3F555E7F9EBEBEE1BB32D8AA00AAA69AE9AE9;
defparam prom_inst_6.INIT_RAM_38 = 256'h082200820AAA0AAA0AA208220AA20AAA0AAA08AA0AAA080272ADFFFFD5552AAA;
defparam prom_inst_6.INIT_RAM_39 = 256'h1D5600001ABE2AAB8AAA028002820A0008000AAA0AA20A000028088208020082;
defparam prom_inst_6.INIT_RAM_3A = 256'hFA18780061B42AA82AAAD5552AAAEAAAAAAB8001E00000005BEAABD60000AAAE;
defparam prom_inst_6.INIT_RAM_3B = 256'h2A00000A8000FFFF80A802A867FEAA6067FFE180387801EE7861E00066000003;
defparam prom_inst_6.INIT_RAM_3C = 256'h1A619F800AAA0000088AEEAA86153554D5552AAD41804180088AAAAAB377AAA0;
defparam prom_inst_6.INIT_RAM_3D = 256'hE7FEB800606061FE1E60060001807FFFFFFEFFFF800067FFFE0006007E607E00;
defparam prom_inst_6.INIT_RAM_3E = 256'hFFF80FFFDFFFFC0FFFBEFFF80FFF85F80660617E01D87F8067F9FFFFC1800001;
defparam prom_inst_6.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80FFFBEFFFB0FFF80FFFBEFFF9CFFF80;

pROM prom_inst_7 (
    .DO({prom_inst_7_dout_w[30:0],prom_inst_7_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_7.READ_MODE = 1'b0;
defparam prom_inst_7.BIT_WIDTH = 1;
defparam prom_inst_7.RESET_MODE = "SYNC";
defparam prom_inst_7.INIT_RAM_00 = 256'hFFFFFF80FFFA6FFFB0FFF80FFFFFFFF80FFFBEFFFA0FFF80FFFBEFFF9CFFF80F;
defparam prom_inst_7.INIT_RAM_01 = 256'h3F3F042909253F21253F3F3F3D253D3F3F2F3F217FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_02 = 256'hAE2AAAFFFFFFFF8001F553EAB8080C002F3C0E1830303F3D192909211806201E;
defparam prom_inst_7.INIT_RAM_03 = 256'hD72CD72A0AAAAAE0607FE07FE000187FE01E0066667FF87FF87FF800002AAFAA;
defparam prom_inst_7.INIT_RAM_04 = 256'hAB2AAAB554D55556AAAAAD2AAD41AAD6AAC1AAAAAAAAAA87FFAAAAAAAAACD72C;
defparam prom_inst_7.INIT_RAM_05 = 256'hAAAAAA01082AA8180001E055535555535554AACAAAC1AACBD4F72AEEAACE152A;
defparam prom_inst_7.INIT_RAM_06 = 256'h0020060000000001FFFFFFFFFFE0002AA02A00000A8000CAAADE405AAAAAAAAA;
defparam prom_inst_7.INIT_RAM_07 = 256'h55FE01F555000076078000781ACAAACAAA80004AAA87FE07FE200627E6200600;
defparam prom_inst_7.INIT_RAM_08 = 256'h552AAAFFFF80007FFF8000007FFFFF800000007FFE7FFE001E00007FFF800075;
defparam prom_inst_7.INIT_RAM_09 = 256'h1F8000001F800099FE00000075755500004E004AAA8000018620067F807FFFD5;
defparam prom_inst_7.INIT_RAM_0A = 256'h8CFFFFFFF083FDDFFFECFCFFFFFFDB1FFFB1FFDF7FFFD9FFF66FDB66DFFFFF80;
defparam prom_inst_7.INIT_RAM_0B = 256'hF80000FCFFFFFBCFF0000C7800FFFFFFFFFFFFFFFF4756DBEC7FEE87FFFFFBFF;
defparam prom_inst_7.INIT_RAM_0C = 256'hFFFFFFFFFF7FFFFFE107FFFFFF5FD780000430FFCF9FFDCFFFF9FF3F9FF3FFFF;
defparam prom_inst_7.INIT_RAM_0D = 256'hFFF7E0201FF7F7F7FF9FB767F8007FFFFFFFFFFFFFFFFF7F7F3FF9FDBA7FC007;
defparam prom_inst_7.INIT_RAM_0E = 256'hFFFFFEAFFC007FEAAFFEFC7FF39FFF01FFFFFFFFFEBFFFFF7FFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_0F = 256'h73E0603FFFFFFFFEBFFFFF7FFFFFFFFFE0605E0605E0605E3FF8FDF77FC007FF;
defparam prom_inst_7.INIT_RAM_10 = 256'hFFFFFFE0605E0605E0605E3FF8FDF77FC007FFFFFEAFD5C0000EAD55FF5F8E06;
defparam prom_inst_7.INIT_RAM_11 = 256'hFFFFFFC03FFFFFFFFFFB7FFFFFFFFFFFFFFFFFFF9FE7F9FEFFC01FFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_12 = 256'h03FFF03FFFFFB7F57FFE03FFF57FFFFBC7F03FFF03FFE27B7FFFFFFFFFE00000;
defparam prom_inst_7.INIT_RAM_13 = 256'hFFD7CFFD40FFD00FFD7CFFD7CFFD00FFDFFFFFFFF17F57FFE03FFF57FFFFBC7F;
defparam prom_inst_7.INIT_RAM_14 = 256'hFE09200FEFFDFEFFDFEFFDFEFFDFEFFDFEFFD00FFD7CFFD60FFD00FFDFEFFD00;
defparam prom_inst_7.INIT_RAM_15 = 256'h0FEAAAC00D7AAAC0000007FFFE7FFFA7FFFE0920000000000007FFFE7FFF87FF;
defparam prom_inst_7.INIT_RAM_16 = 256'hAFAABD5573C00D557028003DC3FCC030C00005EB07EC05EC3DC00FFFF35D3C00;
defparam prom_inst_7.INIT_RAM_17 = 256'hF0000E2B70000E2B70000B0F08FFF3FFC00C03C005D35FAABC7000000D35DFEA;
defparam prom_inst_7.INIT_RAM_18 = 256'hA000003AA0000FAAA000000003FFC0F00AAE20000BFFDAAAF00000000BFFDAAA;
defparam prom_inst_7.INIT_RAM_19 = 256'h5C000FFD5D5703C005FB0D7AA33FC0F0003DCFFFDFEAD555095500000FFAAFAA;
defparam prom_inst_7.INIT_RAM_1A = 256'h400093C005542000AFFFF0000000055C0B0F0000C44409D7AFFFF00005555555;
defparam prom_inst_7.INIT_RAM_1B = 256'h0A070E05CAA55555400000000FCF5AFF5EAE2D54C55509D7AFFFF00035557555;
defparam prom_inst_7.INIT_RAM_1C = 256'h500000808008A02AAFAAAFFFFFFFFAAAA03000003FEB7A57A107C700701D5000;
defparam prom_inst_7.INIT_RAM_1D = 256'h701FF0EABDAF0423F000000000000D7AAFEADAAAA00000000AFD557000000555;
defparam prom_inst_7.INIT_RAM_1E = 256'h0CF5C03DC35F537D5DFAC57ACFD2AAAAAA87FFFD5FD2CFF405555387F57FFDD4;
defparam prom_inst_7.INIT_RAM_1F = 256'hF00080C0F7D5555550C0300FFEB5DEB15A203C000000000000000D6550C3330F;
defparam prom_inst_7.INIT_RAM_20 = 256'hC00F0300C3C0030CC3FFC0FFF0FF7FF00FD70DCFFF00000000000FFF0FD5503F;
defparam prom_inst_7.INIT_RAM_21 = 256'h00000FF000000F0000A00FFF2330C3000300C0F0CFAABDAC00000E40000013FF;
defparam prom_inst_7.INIT_RAM_22 = 256'h200020000A8A002008A2000002ACA00000000FFFF000000000A0000005595004;
defparam prom_inst_7.INIT_RAM_23 = 256'h082A002A08080020008A02080002000800A882220000020020200A20222A0200;
defparam prom_inst_7.INIT_RAM_24 = 256'hE7DF789F5787BEFAEBAF401401440451C5BCA452219200000000882A88002A0A;
defparam prom_inst_7.INIT_RAM_25 = 256'h5A40807C2659E0605A1E240007B6DB6802175FB3EA7AEFDEF7BDEDD87F7DDB7F;
defparam prom_inst_7.INIT_RAM_26 = 256'h90001B6A312D0C3C0DCCC00000302B589555568781B4200081BB991C11046FFF;
defparam prom_inst_7.INIT_RAM_27 = 256'h17C27E7818989A1806F8F03120000000000000000000000883BC625818789BB9;
defparam prom_inst_7.INIT_RAM_28 = 256'hFF7BDEAF44AADAEABD397ABCB95F5EAC95BDF004A46B5B5EDC5EC4B944454A3E;
defparam prom_inst_7.INIT_RAM_29 = 256'hDF0BF1ED989081F4FFFFDF74EA9996997BA5126C48AEBB5B55BDEF7AB6FD4EF2;
defparam prom_inst_7.INIT_RAM_2A = 256'h111111111BA99101328FFF9F5D557EF64DABE6FB7FF7E83D7FBE03DDBF4BF1ED;
defparam prom_inst_7.INIT_RAM_2B = 256'h399D48FF8DD5D1D29DBEB1EAFFBFFFBB5FFE520B2592C964F3CF3CF496EDB55D;
defparam prom_inst_7.INIT_RAM_2C = 256'h554FE53FEAD71BDC844370DECBB79FEB5C1B27FBFCAE56ED32A7FF5D7DA9BFBA;
defparam prom_inst_7.INIT_RAM_2D = 256'h18C6318C610806DA24F51FBCBB527CBEFADBD973F8599A43B96646DA6CD5CF9F;
defparam prom_inst_7.INIT_RAM_2E = 256'h881E703F001FE007C037E042100550150504104445140001441551004500145B;
defparam prom_inst_7.INIT_RAM_2F = 256'h0047026BBD7DAAF17638C11BEF5DC0DC0980702601DF72BF72BA910938C33A81;
defparam prom_inst_7.INIT_RAM_30 = 256'hF5404E402B02C7421D0D0E83D8E09C8C07232B04AB574D676BA7D57D505C00F1;
defparam prom_inst_7.INIT_RAM_31 = 256'h5A533104909108208E08425AC428812AC4358130D55D5354928DC51A9176BF57;
defparam prom_inst_7.INIT_RAM_32 = 256'hD55555400013555D0500000000000003979538B50AD2AAD51C4A806826629608;
defparam prom_inst_7.INIT_RAM_33 = 256'hDAB5AB430202F61A34EEE4BB2200533B20AC30868D3868D0800068D3868D0830;
defparam prom_inst_7.INIT_RAM_34 = 256'h8A548A549B66AD9A49956C000F952A1843E8530202410A4900040015BB76F6DE;
defparam prom_inst_7.INIT_RAM_35 = 256'h0199D77FC020200020002122E9AE89997125DA20489AE980925491220A548A54;
defparam prom_inst_7.INIT_RAM_36 = 256'h08178BC0000743A0840000542A500083E1F0FFAA342A2A2BA8A8003914111410;
defparam prom_inst_7.INIT_RAM_37 = 256'hD76BB08890408028908004041020001400C082118825FF1A8D417C38542A7058;
defparam prom_inst_7.INIT_RAM_38 = 256'h0B1AD016B4E5AD68000024C013686EFBBFCBB0169A0A81561511111111600B2E;
defparam prom_inst_7.INIT_RAM_39 = 256'h1000D6B5AA6B5AD6B5052940028D55400001AD6B401AD6B5AD49014A00147038;
defparam prom_inst_7.INIT_RAM_3A = 256'h009B43D9804D680B5A714B5A28444026D0D104D685AD388804DA1CC03004DA12;
defparam prom_inst_7.INIT_RAM_3B = 256'hAAA9252940028E070184223880098026D0DDD1C3BCEF035AD2AEB4E52D68A111;
defparam prom_inst_7.INIT_RAM_3C = 256'hDE4111044411141415100011138505515540000A00A082AA20007A36555082A8;
defparam prom_inst_7.INIT_RAM_3D = 256'h28088228A8A00A8D9762800365D8A00132AA7115500000000204437775DF75DD;
defparam prom_inst_7.INIT_RAM_3E = 256'h380000297841C0A00DDFF7F5D77E000808B0F50055607F31D32ABED355663E87;
defparam prom_inst_7.INIT_RAM_3F = 256'h002000000000000000D500005511631C0E0320000088100568743A132AA850C4;

pROM prom_inst_8 (
    .DO({prom_inst_8_dout_w[30:0],prom_inst_8_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_8.READ_MODE = 1'b0;
defparam prom_inst_8.BIT_WIDTH = 1;
defparam prom_inst_8.RESET_MODE = "SYNC";
defparam prom_inst_8.INIT_RAM_00 = 256'hFFFFFFFFFD050A89642625948195134245114E842AFAFAFAFFF36CFFFFFFF800;
defparam prom_inst_8.INIT_RAM_01 = 256'h60282A4F0CD904104104820900C102C55F8C444C2840C00002DFF03F10C02004;
defparam prom_inst_8.INIT_RAM_02 = 256'h51023218891239000444CE7281149A4D241A49293187F608236880022C92CD10;
defparam prom_inst_8.INIT_RAM_03 = 256'hB2203080002642482AA0022119884CE75880A01DF75A7D250E2880F77F7D5257;
defparam prom_inst_8.INIT_RAM_04 = 256'h1303898000C622329894412511089A3B0231C0C011B31113953108098C44C4E3;
defparam prom_inst_8.INIT_RAM_05 = 256'h72871550049828B40888A049249A96890110920821390B442E25C11324421420;
defparam prom_inst_8.INIT_RAM_06 = 256'hAA88608010783840155007307020000028F471C089A06094951E6065C40AB632;
defparam prom_inst_8.INIT_RAM_07 = 256'hD2155C211C5168823212045C41501505414E7258A92C8C08A3C454A406240403;
defparam prom_inst_8.INIT_RAM_08 = 256'h8849289001100110999886E48B5113791498C462403F064A202AA40C1B914875;
defparam prom_inst_8.INIT_RAM_09 = 256'hA154A00A0A22720D8898484444003622212F08CE173F940CE44A22221000CD88;
defparam prom_inst_8.INIT_RAM_0A = 256'h732090C70064526C5F7E04584440806C44C20622000B1130841888018B1130B8;
defparam prom_inst_8.INIT_RAM_0B = 256'hE0A1424999513CB16B49411208205AA5C32E2731CD0092912C521782070B6E44;
defparam prom_inst_8.INIT_RAM_0C = 256'hE78C8A42379420A9BCA46681234436591604E6F646C7010D6E48FC71F3F94198;
defparam prom_inst_8.INIT_RAM_0D = 256'h2FD908F74C9500F020C943CA33834A11D33C452809E01158B8446266E315E28C;
defparam prom_inst_8.INIT_RAM_0E = 256'h3893CFD64433C92281E44192079467069423A6788A5413C022B1708A4089238B;
defparam prom_inst_8.INIT_RAM_0F = 256'h619C826A773A92470396DC596E0A888B1090260866442406252B00B3CEA40892;
defparam prom_inst_8.INIT_RAM_10 = 256'hE8BFE8D294C78F921A915369CC739FC12970250F160E1847218A9DCEA499E2C8;
defparam prom_inst_8.INIT_RAM_11 = 256'h109A2858F31622C5848131334E03DC5CC598F3050404DA888E471F681067F742;
defparam prom_inst_8.INIT_RAM_12 = 256'hFFE1364C4D4B49B9A889328421133CA18B322944828F02169A69882C164F342C;
defparam prom_inst_8.INIT_RAM_13 = 256'h4466B004CA108C72862CC9A5368A1C085913608C51429899C48F00E0884D0036;
defparam prom_inst_8.INIT_RAM_14 = 256'hD9DAF9691F5401084B21AF7F2076213CB9FEC38220600094CFFEFC1001309464;
defparam prom_inst_8.INIT_RAM_15 = 256'h98E29B44110409908D82673299386260C6A33D897E3DDB77018564698EEF87CC;
defparam prom_inst_8.INIT_RAM_16 = 256'hC0991A37788975C2931C53688220864C85036099C8A45CC9C11011BBC44BAE16;
defparam prom_inst_8.INIT_RAM_17 = 256'h4E267AA432891E1BE0C7247879C800834A126253F038DBC4BAE1491E29B44110;
defparam prom_inst_8.INIT_RAM_18 = 256'h80774822CA03042828660480CD4590D922426CC7C052A34E0F0143FF1F23C82D;
defparam prom_inst_8.INIT_RAM_19 = 256'h997444D1C1B1D73F183045D9474C18228CF46D5002A2AC9C98C636DBCD8A5004;
defparam prom_inst_8.INIT_RAM_1A = 256'hB3B91D0392DC14DCD9A000121C4907722930C87A9B118904D99F3B02D9AA9030;
defparam prom_inst_8.INIT_RAM_1B = 256'h21A2C0248003136C48927A1B58A26288EC84F000000000000CD26AC1600070D5;
defparam prom_inst_8.INIT_RAM_1C = 256'h39544105A8EF208C1064EEF006289149BCC0950798804CD096660181A4523892;
defparam prom_inst_8.INIT_RAM_1D = 256'hE4E3478620A0421148AA90948800C000CE410460082C0603010820467A642042;
defparam prom_inst_8.INIT_RAM_1E = 256'h1950810C90A2A10214220FCAD21E6811585488CE4DD4305A495A13983330A2CC;
defparam prom_inst_8.INIT_RAM_1F = 256'h0461280611A20429A0606860145A19A5033A173968B70C618CE6618884494A2A;
defparam prom_inst_8.INIT_RAM_20 = 256'hF834DA8891088422C4E146C1970623080C82B4A4D8BEFC08C8E81AC8855B6426;
defparam prom_inst_8.INIT_RAM_21 = 256'h76E63227664D821148A406EBBBBE236E0999997F448408C9D080F416470F32C8;
defparam prom_inst_8.INIT_RAM_22 = 256'h85030A06140C28185030A061500054089C6926145A4A3847091B5046046E3811;
defparam prom_inst_8.INIT_RAM_23 = 256'h1F1A780900C0D280C68540634018D030A06140C28185030A06140C2A336C8241;
defparam prom_inst_8.INIT_RAM_24 = 256'h808475896F862090C0B2C30C29171D177057AF15D3C689168A4D804550623335;
defparam prom_inst_8.INIT_RAM_25 = 256'h010205B71244C5BC240A208E91000D414412211B1160C08B0051122281849028;
defparam prom_inst_8.INIT_RAM_26 = 256'h0010020821C7404379D32808444009880102CEA8042012240608A84180035008;
defparam prom_inst_8.INIT_RAM_27 = 256'hCD2CA018002DE29003800B65A8C61861060C61061020010C1046106006184182;
defparam prom_inst_8.INIT_RAM_28 = 256'h000001E8000003E000000B0000003E002800FC0030006C0038926D8309CD2380;
defparam prom_inst_8.INIT_RAM_29 = 256'h9E493578C8285555534154401A00018004C0000B000500002002DE000000003C;
defparam prom_inst_8.INIT_RAM_2A = 256'hA4B7684CF2B76DB60CD4988B6DCCDAA8B1F18491A24244848051EE09CA3F5B9A;
defparam prom_inst_8.INIT_RAM_2B = 256'h005500F055F0A055200550055005500550055004255596DC64A7BD305CCF7A64;
defparam prom_inst_8.INIT_RAM_2C = 256'hEFECCDDCCDCCCD110000111101109898989898989889898989898989AFA50055;
defparam prom_inst_8.INIT_RAM_2D = 256'hEBBBB43FE9BBF477D767EB8FFAEE7D8BFA777EA3FEFEEFFEFFEEFFEEFFEEEFFE;
defparam prom_inst_8.INIT_RAM_2E = 256'hFA37EB9DF49FFAE77D27FEB37E9CFFACDFA73FE99FFA67FE99FFA67FEBBBB43F;
defparam prom_inst_8.INIT_RAM_2F = 256'hC2C4A65E63A7CE97FFB07BD5C289733E4755555555550AA954AA5677EB1FF5CD;
defparam prom_inst_8.INIT_RAM_30 = 256'hCC89DFE01E181D7FFFDFBFFFEBF4BA5FFFF0E1D57871E3CF9F4F9D2FFF63DBD5;
defparam prom_inst_8.INIT_RAM_31 = 256'hB10A00AA014141EBEB41413C7492FFAFFF492EB8751400BC7A3D145028BAF88C;
defparam prom_inst_8.INIT_RAM_32 = 256'h2AAA80FF9C3FABFFFFFFFFFFFFFFFFE47FFFFFFF91FFFFFFEB041EBEB4141EBE;
defparam prom_inst_8.INIT_RAM_33 = 256'h80007FFF807828787FF8114451FFD1FFFFE411E47FFFFFFFFFA07E967FEA8000;
defparam prom_inst_8.INIT_RAM_34 = 256'h7FFF9AAA9AAA9ABE1AAE9AAAFAAAAAAAABAAABAA9EAAAAAAAAAE0780078287FF;
defparam prom_inst_8.INIT_RAM_35 = 256'h2AAE07E007881155115501FF80007FFF81F802787FE0000011FFFFE47FE40000;
defparam prom_inst_8.INIT_RAM_36 = 256'hAFFA88020822008200A01AAAFAAA9D561D561D567FFF9AAA80001AAA9AAE9ABE;
defparam prom_inst_8.INIT_RAM_37 = 256'hECABEAABEACCACAB72A9F61DEEA3F555E7F9EBEBEE1BAAAB8AA00AAA7FAFFAFF;
defparam prom_inst_8.INIT_RAM_38 = 256'h08220082088208220A8208220822020208220A820AAA08026B2BFFFFD5552AAA;
defparam prom_inst_8.INIT_RAM_39 = 256'h1D5600001ABE2BAB880200A00082080008000AAA0822080000A0080208020082;
defparam prom_inst_8.INIT_RAM_3A = 256'h18E007E0183028002AAAD5552AAAEAAAAAAB8001E00000007AFAEFD60000AAAE;
defparam prom_inst_8.INIT_RAM_3B = 256'h2A0000028000FFFF80A000A00001546000001E005619E7AE07E1980061EC1F82;
defparam prom_inst_8.INIT_RAM_3C = 256'h789E00000AAA8000088AEF2A81812AAAD5502AB506000600088AAAAAB377AA80;
defparam prom_inst_8.INIT_RAM_3D = 256'h8006DE003F807E6299FFE60006007FFEFFFEFFFF800000007580780075800000;
defparam prom_inst_8.INIT_RAM_3E = 256'h8017E80100801008011A8017F8011CF807E0673E01D81D8000007FFFBE000001;
defparam prom_inst_8.INIT_RAM_3F = 256'h017E801428014280142801428017E8017F801418016F80100801418016B8017F;

pROM prom_inst_9 (
    .DO({prom_inst_9_dout_w[30:0],prom_inst_9_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_9.READ_MODE = 1'b0;
defparam prom_inst_9.BIT_WIDTH = 1;
defparam prom_inst_9.RESET_MODE = "SYNC";
defparam prom_inst_9.INIT_RAM_00 = 256'h17E8017F801418016F8017F801008017F801418015F80100801418016B8017F8;
defparam prom_inst_9.INIT_RAM_01 = 256'h213F042109252121250929253925251125393F217E8014280142801428014280;
defparam prom_inst_9.INIT_RAM_02 = 256'hAFABAAFFFFFFFF800075539AAE140C003D3C0C0C20203F25092109210C0C200C;
defparam prom_inst_9.INIT_RAM_03 = 256'hD72CD72A0AAA8AFFE01F8000007FFE7FE001E06666619866187FF800002AAE2A;
defparam prom_inst_9.INIT_RAM_04 = 256'h52AAAAAAAAD55035AAAAAAAAB506AAB5AA86AAAAAAAAAA87FFAAAAAAAAACD72C;
defparam prom_inst_9.INIT_RAM_05 = 256'hAAAAA801082AAA1FFE07F8552CD554D3552AAAD2AA86AACF4AF7556F2AD38155;
defparam prom_inst_9.INIT_RAM_06 = 256'h0020067FFF8000781FFFFFFFFFF8002A802A0000028000DAAADE404AAAAAAAAA;
defparam prom_inst_9.INIT_RAM_07 = 256'h5577E07555000075E780005E07EAAACAAA80004AAA801800062006207E200600;
defparam prom_inst_9.INIT_RAM_08 = 256'h552AAAFFFF8000755500000007CAAA8000000020062006006600007FFF800075;
defparam prom_inst_9.INIT_RAM_09 = 256'h0780000007800099FE7E00001D7555007FD8004AAAFFFE006620067E007FFFD5;
defparam prom_inst_9.INIT_RAM_0A = 256'hFB0000003F7C009601EB8100000015E018CCC0225803D70319BD7C0938000000;
defparam prom_inst_9.INIT_RAM_0B = 256'hF00000C0800DFC70DFC70F8470FFFFF80000000007F2082F93C3997E000000D5;
defparam prom_inst_9.INIT_RAM_0C = 256'h00000000000000007EF83F8FE2388E000001CF00006101000000101090403FFF;
defparam prom_inst_9.INIT_RAM_0D = 256'h38FE1FDFE1FCFE1BDF6054F807FF80000000000000001FCFE1DDF602A5803FF8;
defparam prom_inst_9.INIT_RAM_0E = 256'h0000355803FF80355803D7800D6000FE00000000028000000000000000000001;
defparam prom_inst_9.INIT_RAM_0F = 256'hAC1F9FC00000000280000000000000002000120001200013DFF702D7803FF800;
defparam prom_inst_9.INIT_RAM_10 = 256'h0000002000120001200013DFF702D7803FF80000035EAB3FFFF35EAB25FAF1F9;
defparam prom_inst_9.INIT_RAM_11 = 256'h00000FC03F00040FFFF7C1101C01E020087A1E87E7F80601003FE00000000000;
defparam prom_inst_9.INIT_RAM_12 = 256'hFC000FC00000E81AC001FC481AC4812C780FC000FC001F6E8000000000000000;
defparam prom_inst_9.INIT_RAM_13 = 256'h00283002BF002010028300283002FF00200000000F81AC001FC481AC4812C780;
defparam prom_inst_9.INIT_RAM_14 = 256'h7E00000FD00285002850028500285002FD002FF00283002DF002FF00201002FF;
defparam prom_inst_9.INIT_RAM_15 = 256'h0FEAAAC00D7FFAC0000000003E000560007E00000FFFFF000000003E0006E000;
defparam prom_inst_9.INIT_RAM_16 = 256'hAFAABF5DF0000F5DF0000CF5C30CC030C00005FB09AC35EC0CC00FFFFF5FFC00;
defparam prom_inst_9.INIT_RAM_17 = 256'hD0000BFF50000BFF50000FC330FFF3FFC00C0C7005FF5FAAB3C000000FF5FFEA;
defparam prom_inst_9.INIT_RAM_18 = 256'hA000003AA0000FFAA000000003FFC03C0FFBF0000AAAFBFFD00000000AAAFBFF;
defparam prom_inst_9.INIT_RAM_19 = 256'h00000AFD5355C3000A6B0D7FF33FC03C0CF5CFEAAFFFDA550AA500000FAAAFFA;
defparam prom_inst_9.INIT_RAM_1A = 256'h30002C7005502401AAAAA0000000055C0FC3300034440957A0808C000AAAA000;
defparam prom_inst_9.INIT_RAM_1B = 256'h0857045700295A95500000000AFF5FCF5EBFF555C5550957AAA08000DAAA9000;
defparam prom_inst_9.INIT_RAM_1C = 256'hA0000AAAA00A200AAFFAAFEAAAAAAFFBFFC000003FEB7A57A51734417407F3C0;
defparam prom_inst_9.INIT_RAM_1D = 256'h757FF0EBD7ECC3FC0000000000000D7FFFFFDFFBF00005555FFD557000000AAA;
defparam prom_inst_9.INIT_RAM_1E = 256'h303DCCF5C37D535F557ACDFACFD000000007FFF40FD2CFFD50000387F01FFDD4;
defparam prom_inst_9.INIT_RAM_1F = 256'h0AAA00C03AAAA3C000C0FF357D77AC20C00AA0000000000000000D60030F00C3;
defparam prom_inst_9.INIT_RAM_20 = 256'hC03C0300C300030CC300C0FFF0D55FFC05570F000000000000000555C57FFFC0;
defparam prom_inst_9.INIT_RAM_21 = 256'h000000A0000005F00A000FFF0300C3000300C030CFFFD7EC0FF00E4000001030;
defparam prom_inst_9.INIT_RAM_22 = 256'h4442244014820080002000000555455540000080800000000AA000000AAA9004;
defparam prom_inst_9.INIT_RAM_23 = 256'h44000000542A02854000004C4414220846A20482000020000022D486002A2684;
defparam prom_inst_9.INIT_RAM_24 = 256'h4B69019E47A8104104110015101151107C208347D803000000008C0044442828;
defparam prom_inst_9.INIT_RAM_25 = 256'h9E20002D334010509E01244231A69A788FB311F39AD2DA14A5ADB4056DA40012;
defparam prom_inst_9.INIT_RAM_26 = 256'h0004524C614914024810500AA428210826666780410718CE41002012082E4319;
defparam prom_inst_9.INIT_RAM_27 = 256'h128238043410921210B809687800D556BBFFFC01FE044C4D4104CA9228041002;
defparam prom_inst_9.INIT_RAM_28 = 256'hDA52D6B1770894DD8B91A338D1956AC859D40294A4129E10F78CB75DE0859A42;
defparam prom_inst_9.INIT_RAM_29 = 256'hE2432161AA1494E4E69B6904C4614A003D200244991763FDFFC94A5ADB2D8840;
defparam prom_inst_9.INIT_RAM_2A = 256'h222222331B3BB10203CFFF1A1E877078AA33F4AD99999814524A4D8802032141;
defparam prom_inst_9.INIT_RAM_2B = 256'hA19148CBCF413FAEFA90B815014284910D32172160F8583E14714718BB02C992;
defparam prom_inst_9.INIT_RAM_2C = 256'h66D8042F48F309E2ACA78119893D08426D0330C2050364C067A8500439190080;
defparam prom_inst_9.INIT_RAM_2D = 256'hCE739CE73A42069C3C46047CABC3E030C37D1131503B395E3EC0CC1349101210;
defparam prom_inst_9.INIT_RAM_2E = 256'h118EFB9551FE015991DFE6409005554005501505041044451400014415510041;
defparam prom_inst_9.INIT_RAM_2F = 256'hFCF81D0BE1D42AC1D8280102A87780617C2E8172AF1542FC75272312F1163503;
defparam prom_inst_9.INIT_RAM_30 = 256'h5F616E5536FAD0AB42EDB00800126583DD65F30424C101E12082822820EFAE7E;
defparam prom_inst_9.INIT_RAM_31 = 256'h00530100104008378178C080116A0040100021BBFFEFABA862576AAEC5DE55F5;
defparam prom_inst_9.INIT_RAM_32 = 256'hEBEBEFEFFFFBABBEAE000000AAAAAAA085108D95E050005504D1481466401608;
defparam prom_inst_9.INIT_RAM_33 = 256'h000000010202B4DBB4291D3B2208DFFB2001D0B6ED0B6ED180036ED0B6ED08BF;
defparam prom_inst_9.INIT_RAM_34 = 256'h803018301356ED5A002002D5AD952A1843085502020AD2258836209000000801;
defparam prom_inst_9.INIT_RAM_35 = 256'h21805D556A8AAAAA8AAA8303F7D7400012311330C0FF7DD8D37691221B768036;
defparam prom_inst_9.INIT_RAM_36 = 256'h020F87CBEA85E2F192C550D46A500007E3F0FFFDFDF5F5D5D950000CEA31143B;
defparam prom_inst_9.INIT_RAM_37 = 256'h000BB020216030289000040458000020002002000020AA000000541040201000;
defparam prom_inst_9.INIT_RAM_38 = 256'h001AD2C6B425A00006B46836AF68EEFFFB8EE156308AB156100000000016BB00;
defparam prom_inst_9.INIT_RAM_39 = 256'h00000000026B5AD6B548421084000000000000000B5AD6B5AD70421084200000;
defparam prom_inst_9.INIT_RAM_3A = 256'hB57B4351002D6AD35A10200140452D5ED0F982D699AD08A5ABDA18800DABDA12;
defparam prom_inst_9.INIT_RAM_3B = 256'hAAA96842108400000004C23800906D5ED1FD79600000023AD276B42080050314;
defparam prom_inst_9.INIT_RAM_3C = 256'h5C00000000000540140000400080055155400018AA0080000AA8EE2000000002;
defparam prom_inst_9.INIT_RAM_3D = 256'h02AAA8800200000FE6602AA3F99A0AA8233215555000000003804377F77775DF;
defparam prom_inst_9.INIT_RAM_3E = 256'h0800002D7BF5FA1D0FF777FD5FF600000A803560C460FB211BB3371BE608B703;
defparam prom_inst_9.INIT_RAM_3F = 256'h000200000000000AD67700000005481C0E02BBB8000025ED6875FA000000AFBB;

pROM prom_inst_10 (
    .DO({prom_inst_10_dout_w[30:0],prom_inst_10_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_10.READ_MODE = 1'b0;
defparam prom_inst_10.BIT_WIDTH = 1;
defparam prom_inst_10.RESET_MODE = "SYNC";
defparam prom_inst_10.INIT_RAM_00 = 256'hFFFFFFFFFD6528AB54AEAD529AB1755A57D46B1518FEFEFAFFFC82FFFFFFF800;
defparam prom_inst_10.INIT_RAM_01 = 256'hF9E7B9AAC8C26D26DB4936934CD56EB65D6E775EAD708000000F05F0C00020E0;
defparam prom_inst_10.INIT_RAM_02 = 256'h270FBADDB9C2B9655D7D5F74CF969F4FB4CF683D1DD7F7AAEBAAABAF6ED074B5;
defparam prom_inst_10.INIT_RAM_03 = 256'hDA465A871C77CC91DD5F9AED7FBBFD76A1184DA2A88A0A8800A2AA8AAA8002A2;
defparam prom_inst_10.INIT_RAM_04 = 256'h75ADD9B57FF7AAEE9EC332267D6AA8F75EF28C36DDDFF55757FFFDAB95D7F55A;
defparam prom_inst_10.INIT_RAM_05 = 256'hEEBF6AAADC51EA953BBBEFFFFFF797BAE7D67FFBEFE77BDDAC47ED5745587AD4;
defparam prom_inst_10.INIT_RAM_06 = 256'h5578231502A15DC2EAAAD4630DB51125EA959682AAAD5316B56AED5D4889801D;
defparam prom_inst_10.INIT_RAM_07 = 256'hA2A36F60DD415BB9BD06DF55279EB49E7B75A3D69A3741BEBEB7D654567CDCCD;
defparam prom_inst_10.INIT_RAM_08 = 256'hBB016BDD5C491802EABA0DBC38DE9AE743B143D8B3A43A91555D53C04618CA7C;
defparam prom_inst_10.INIT_RAM_09 = 256'h85DF999ABABBBA35EABB03755161D7AAEC09BAC9AAC8C816C1EF9BAAC30835EA;
defparam prom_inst_10.INIT_RAM_0A = 256'hAC48565547F57FFDB5BEA57A646891EF5558D7AAB27BD556335EAAC07BD55622;
defparam prom_inst_10.INIT_RAM_0B = 256'hAC3507EED74D2C815BFCEB865025D55BEEB9BAFBB44DA601F73A5ED647AFBC65;
defparam prom_inst_10.INIT_RAM_0C = 256'hAEAEB9BB80C80D460640B330D514D9DED8375DD035FD255F5DEB657850AF32BF;
defparam prom_inst_10.INIT_RAM_0D = 256'h6F556EBEDE3F2B77E7594EBABA2E8CD54D2B7F2B7EA0C7726BDCBFABBD17AE6B;
defparam prom_inst_10.INIT_RAM_0E = 256'hAFDBDBF574BADC7656EBCEB29D75745D19AA9A56FE52FD41CEC4D7BADEB99AFB;
defparam prom_inst_10.INIT_RAM_0F = 256'h3F6A7ABA42568D5A1FFFF9FFFCFB8384660F33032662000627929BAAABACEB99;
defparam prom_inst_10.INIT_RAM_10 = 256'hEFFFEDC5CA146E4D596D12092FBDECAC1CFC5C1409B50FDA9EAE9095A35E8034;
defparam prom_inst_10.INIT_RAM_11 = 256'hF7FBA5C84D09E018F078DFF5CA0EFB7942680D2D2D55AEB6B555572AE1F7B77F;
defparam prom_inst_10.INIT_RAM_12 = 256'h77EFF2DB75152D4C0EBB3675EF555D9D791BB976EA773BF269A2A3A4F0FFF3E4;
defparam prom_inst_10.INIT_RAM_13 = 256'h5DAB36CCD9D7BDF675E46FE5DB29FCEFC3DF27BFDD2E6FFAFC9D0627BB566CF7;
defparam prom_inst_10.INIT_RAM_14 = 256'h6EEC6B01144DDC442350AF249815AD518AE08088461B2BD6117EFC00033BB237;
defparam prom_inst_10.INIT_RAM_15 = 256'h046A0ADDCDC731A8341BAA060508842CB4DD5D6B25B9B86ECC266A07A88EB677;
defparam prom_inst_10.INIT_RAM_16 = 256'h731A81C280A236F6408D415BB9B8E38D40ED06EA8581402846232D415051B7B0;
defparam prom_inst_10.INIT_RAM_17 = 256'h6230CBB16780F2C32D1503CB054D8CE9E445AE4A4836C1051B7B2046A0ADDCDC;
defparam prom_inst_10.INIT_RAM_18 = 256'h378697156444DDB353B0E11E029809FA5AB6CE0E42A11662392E88D8C195033F;
defparam prom_inst_10.INIT_RAM_19 = 256'hA3514D9715AD43E754FB5F9F35DA7DAFB5758408C66EE495A575E4831E6B3B0D;
defparam prom_inst_10.INIT_RAM_1A = 256'h04A97B754640F3B6BFBE490ACA5ADF4E8763BDF7F50F62DF4BAF723C43754F3A;
defparam prom_inst_10.INIT_RAM_1B = 256'h94821369800E1F815FD7E8DF3BEAF8ABDEA4C4D4A15A84626139DBA008000FCB;
defparam prom_inst_10.INIT_RAM_1C = 256'hA18B90940D201AD40FB5DD56AAEBD70DD6FBB6F2D1212E3A80B4F7AD45C2B50A;
defparam prom_inst_10.INIT_RAM_1D = 256'h1847DA8C4405DA57656CC5391C98EC76BE9097763040601018EC85DABAB7845B;
defparam prom_inst_10.INIT_RAM_1E = 256'h05607686949B9A4DF308427B20639ED750BCE776EFEE02EECEB0FD763982AAE0;
defparam prom_inst_10.INIT_RAM_1F = 256'h4C059D283DB0986B062626219DDAC2728FDED529CB7518A311CBED6BB55180AD;
defparam prom_inst_10.INIT_RAM_20 = 256'h28487A79593BA4E55CA8DAF5DBF5FDF9EEB2587FFB6B7D4B2F795DD6BDCFB4B3;
defparam prom_inst_10.INIT_RAM_21 = 256'h599B14E5193B8351A8D4677FD8D73AED3F5427C9E9E0576942A62D53772FB24F;
defparam prom_inst_10.INIT_RAM_22 = 256'h67604EC99D813B267604EC99DA5B6699636CF126A48EE439BF228F75B55BCD35;
defparam prom_inst_10.INIT_RAM_23 = 256'h10BA42BDF812767933B73C09D3267604EC99D813B267604EC99D8139BD26AF72;
defparam prom_inst_10.INIT_RAM_24 = 256'h77A37CAB2CAF10F4CBF9825EA4D9BD3ED993B53661F6BB26B9F4A3D54B5BEDF7;
defparam prom_inst_10.INIT_RAM_25 = 256'h51168FEE524AAAAEB39DF84A58F73F73BF08E8D9D7F966CEE5CD93AFF2DC9339;
defparam prom_inst_10.INIT_RAM_26 = 256'h1C71861060C3404225994C855D50AAAA156A1AED1EC6D264FC36E685D562C3ED;
defparam prom_inst_10.INIT_RAM_27 = 256'h13910B00CA3C108B01F28F17B8741015841000010400030C30471C71C75C71D7;
defparam prom_inst_10.INIT_RAM_28 = 256'h7FC3BE05FF8EF817FE3BE05FFCEF81FF87FE01FFCFFF83FFC6F775CF6E139746;
defparam prom_inst_10.INIT_RAM_29 = 256'h8F221519DBAB5555554D55FFE0FFFE7FF03FFFF0FFF0FFFFF7F821FFFFF7FFC1;
defparam prom_inst_10.INIT_RAM_2A = 256'h85F8375DEB489240EE30671A16ABB6FADD9DBA75ABF7D7EC71D81F0CE01B7E0A;
defparam prom_inst_10.INIT_RAM_2B = 256'hFFAAAAFAFFFFFFAAAAAFFFFAAAAFFFFAAAAFFFF96F54DB4DB6D09C1640A1382C;
defparam prom_inst_10.INIT_RAM_2C = 256'hFEEFFEEEEFFEEF3333332222ABBBFFEEEEFFEEFFEEFEEFFEEFFEEFFEAAAAAAFF;
defparam prom_inst_10.INIT_RAM_2D = 256'hFBBBBC3FF9BBFC77F767FB8FFEEE7F8BFE777FA3FFEEEFFFEEEEFFFFEEEEEFFF;
defparam prom_inst_10.INIT_RAM_2E = 256'hFE37FB9DFC9FFEE77F27FFB37F9CFFECDFE73FF99FFE67FF99FFE67FFBBBBC3F;
defparam prom_inst_10.INIT_RAM_2F = 256'hFC35F87796E5CA95FEFF83DFFC6BFC6FAD5555555555C6954AA55677FB1FFDCD;
defparam prom_inst_10.INIT_RAM_30 = 256'hCCCFBA1E01F81F4EFDEEFD7FBD54AA57EFDFBF7FEFDEBD72E5CB952BFDED93DF;
defparam prom_inst_10.INIT_RAM_31 = 256'h000AAA0001540000000001D75FFFA924AA4924AFDFFFFFFF8FC71C7FFFFBECC8;
defparam prom_inst_10.INIT_RAM_32 = 256'h7FFFC83F9C3FFFFF80007FFFFFF87FE47FFF87FF91FFFFFF80000AAAAAAAA000;
defparam prom_inst_10.INIT_RAM_33 = 256'h80007FFF807868787FF81144000051FFFFE411E407F87FFFFE837E967FFFD555;
defparam prom_inst_10.INIT_RAM_34 = 256'h2AAA9AAA9AAB9EBE1AAA9AAEAAAAFFFFAAAAEAAA9EAAAAAAABAE0780078287FF;
defparam prom_inst_10.INIT_RAM_35 = 256'h2BAE0782878811501155007FAAAAFFFFA87802787F80006011FF87E47FE40000;
defparam prom_inst_10.INIT_RAM_36 = 256'hA6BA0AAA0AAA008200A01BABAAAA9D561D561D562AAA9AEA80001AAB9AAA9EBE;
defparam prom_inst_10.INIT_RAM_37 = 256'hEACDECADF2AACACAF2A9F7FDEE03F555E7F9EAABEFFBB2B3802A00026BA6BA6B;
defparam prom_inst_10.INIT_RAM_38 = 256'h0AAA0AAA088208220A020AAA082A020A08220A8208080AAA72B3FFFFD5552AAA;
defparam prom_inst_10.INIT_RAM_39 = 256'h1D5600001EBE2AAB880200280AAA02000AAA0802082A080000280AAA0AAA0AAA;
defparam prom_inst_10.INIT_RAM_3A = 256'h9F805618078000002AAAD5550000600000018001E00000007FABFF580000ABAE;
defparam prom_inst_10.INIT_RAM_3B = 256'h2A8000008002FFFF82880AAA000051800000000059FFFEB8786197E0186D1A61;
defparam prom_inst_10.INIT_RAM_3C = 256'h7A1B80000AAA0000088AEF4A80782AAA80002AD478001800088AAAAAB377AA00;
defparam prom_inst_10.INIT_RAM_3D = 256'h8006D9802E0079FF80007F8061807EBEFEBEFE6067FF80007760000077600000;
defparam prom_inst_10.INIT_RAM_3E = 256'hFFFFEFFFDFFFFC1FFF80FFFFFFFF9CF8786066BE01D81D8000007E602E0067FF;
defparam prom_inst_10.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC1FFF80FFFFFFFFC1FFFFF;

pROM prom_inst_11 (
    .DO({prom_inst_11_dout_w[30:0],prom_inst_11_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_11.READ_MODE = 1'b0;
defparam prom_inst_11.BIT_WIDTH = 1;
defparam prom_inst_11.RESET_MODE = "SYNC";
defparam prom_inst_11.INIT_RAM_00 = 256'hFFFFFFFFFFFE7FFFC1FFFFFFFF81FFFFFFFFFFFFFE1FFF80FFFFFFFFC1FFFFFF;
defparam prom_inst_11.INIT_RAM_01 = 256'h3821043F3F3F213F3F092925313F27132539223F7FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_02 = 256'hAAAAAAFFFFFFFF8001F5538686220C3039071A18102001273F3F3F3F06063F3F;
defparam prom_inst_11.INIT_RAM_03 = 256'hD72CD72AAAAAAA9F80000067807FFE0000001E67E661986618606000002AAE2A;
defparam prom_inst_11.INIT_RAM_04 = 256'h54D4AAAAAA80002D6AAAAAAAD47AAAAB6A9AAAAAAAAAAA87FFFEAAAAAAFED72C;
defparam prom_inst_11.INIT_RAM_05 = 256'hFFAAA001087FFF9FFE1FFE4AAAD2AAD3552AAACAAA9ACAFF2D77556F4AD2F855;
defparam prom_inst_11.INIT_RAM_06 = 256'h0020067FFF81FFFE07FFFFFFFFFE002A002A8000008002DEAADE407FFFAAAAFF;
defparam prom_inst_11.INIT_RAM_07 = 256'h55757875550000755F00004F801EAACAAA81FFCAAA8060000660062018200678;
defparam prom_inst_11.INIT_RAM_08 = 256'h552AAAFFFF80007555000000004AAA8000000078062006078600007FFFE00075;
defparam prom_inst_11.INIT_RAM_09 = 256'h001F80000000009F86780000077555001FE0004AAAFFFE001E200678007FFFD5;
defparam prom_inst_11.INIT_RAM_0A = 256'h047FFFFFFFFFFE21FC1021FFFFFFE01FE4023F8887F8207C8040810C47FFFF9E;
defparam prom_inst_11.INIT_RAM_0B = 256'hF7FFFF3FA493FA093F8003F80000000000007FFFF809A340440C0201FFFFFC02;
defparam prom_inst_11.INIT_RAM_0C = 256'h3FFFF000007FFFFFFFFFC0701C8721800000000000010100000010D0904C3FFF;
defparam prom_inst_11.INIT_RAM_0D = 256'hC73D3FFFF23F3D2420938A07380073FFFF3FFFF3020323F3D222093C5073C007;
defparam prom_inst_11.INIT_RAM_0E = 256'hAAF3CAA73FFFF3CAA73C2873F01F3F01F3FFFF3FF9500000000003FFFF302032;
defparam prom_inst_11.INIT_RAM_0F = 256'h03206033FFFF3FF950000000000200051FFFC1FFFC1FFFC0200C3C0873C0073E;
defparam prom_inst_11.INIT_RAM_10 = 256'h0200051FFFC1FFFC1FFFC0200C3C0873C0072AD550A1543FFFF0A1541A850206;
defparam prom_inst_11.INIT_RAM_11 = 256'hFFFFF7000001F80FFFFDFEFFFFFFFFDFF7FDFF7F9FE7F9FEFF80000000000000;
defparam prom_inst_11.INIT_RAM_12 = 256'h03FE703FE75706653CE7FFB6653B66D786703FE703FE609067FFFE0000000000;
defparam prom_inst_11.INIT_RAM_13 = 256'hFFEFFFFEC3FFE01FFEFFFFEFFFFEFFFFE0000075706653CE7FFB6653B66D7867;
defparam prom_inst_11.INIT_RAM_14 = 256'hC000000FFFFEFFFFEFFFFEFFFFEFFFFEFFFFEFFFFEFFFFE83FFEFFFFE03FFEFF;
defparam prom_inst_11.INIT_RAM_15 = 256'h0FAAAB000D703B00000000003E36DFE36DC00000000000000000003E36DFE36D;
defparam prom_inst_11.INIT_RAM_16 = 256'hBFAAA57FE000057FE0000FD7030FC3FFCF000F3C0DAB05F003000FFFF74D7000;
defparam prom_inst_11.INIT_RAM_17 = 256'hF0000F55F0000F55F00005FFF8FFF000C00C03CC04D747FAC00000000D74D7FE;
defparam prom_inst_11.INIT_RAM_18 = 256'hA000003AA0000FCFA00000000300C0F00F0FD0000AABFF55F0000003FAABFF55;
defparam prom_inst_11.INIT_RAM_19 = 256'h00000FF550D0C0C00F6ACD700000000F0FD70FAA2F00DA550AA500000FAAAFCF;
defparam prom_inst_11.INIT_RAM_1A = 256'hC00003CC0956A556AAAAA00000000570057FF000044409D7A2222FFFF5555000;
defparam prom_inst_11.INIT_RAM_1B = 256'h0C7C0D5C000AAAA9500000000FFD55FFFEB03FFFC55509D7AAA22FFF45556FFF;
defparam prom_inst_11.INIT_RAM_1C = 256'hA00000000008A0002FCFBFAA2AAAAF0FD00000003FEB7A57A7DC0945ED174C30;
defparam prom_inst_11.INIT_RAM_1D = 256'h7FFFF0EB3570CC000000000030000D700F003C3F50000FFFF7FFD5C000000EAA;
defparam prom_inst_11.INIT_RAM_1E = 256'hF03D7FD70D7F50F5703EBFEB0FD255555587FFD06FD2CFFFFAAAA387F907FDC0;
defparam prom_inst_11.INIT_RAM_1F = 256'h000000C0055553C00CC3CED5BEFB5DA0C000000000000000000003FFF33FF03F;
defparam prom_inst_11.INIT_RAM_20 = 256'hC00F03FFC30003FFC300C0D550D5555F055C00000000000000000000B555F000;
defparam prom_inst_11.INIT_RAM_21 = 256'hA00002200000095C00000FFF23FFC3FFC3FFC3FFCF305CF00FF00E4000001030;
defparam prom_inst_11.INIT_RAM_22 = 256'h002080000000000640060000055550000000022220000000000000000AAAA00A;
defparam prom_inst_11.INIT_RAM_23 = 256'h0000446080204420245400000000840200000004440008444408000044000020;
defparam prom_inst_11.INIT_RAM_24 = 256'h91B6EFEF55CBEAFEAFEBFFEAFAABBFFB00000000000000000000080000000020;
defparam prom_inst_11.INIT_RAM_25 = 256'h5DEEC222AABB37675DB354C611659659995DFFD8F7A77CF19C66DBC4B6DBE9B6;
defparam prom_inst_11.INIT_RAM_26 = 256'h402A56D82E9A9366AA22654660B294A54555576CD54318CEDD444454F3CB5155;
defparam prom_inst_11.INIT_RAM_27 = 256'h723BAECD5D76F7751DAD9AFAE7FFCCCD3FFFFC0001EC8409D7485D3726CDD444;
defparam prom_inst_11.INIT_RAM_28 = 256'hB8CE335CF32A9BAAAECEFDA77EDABD6EAD7B398C6223971CBBE53F57B2EEC965;
defparam prom_inst_11.INIT_RAM_29 = 256'h4EACEB1645EAEAB7CB65B6E6DC3BF3A0A6332000000EEF02235319C56DE6F5BA;
defparam prom_inst_11.INIT_RAM_2A = 256'hBBBBBBBB203329919DF63B786E1B383EFFBADF66EEEEF7BEB699EFB6CEECEF16;
defparam prom_inst_11.INIT_RAM_2B = 256'h6979AAD9ABA161479532EFFFD3264D66E6CF54880C4E27018228A0840DE12017;
defparam prom_inst_11.INIT_RAM_2C = 256'h4007D7662EBC6D9512CA555E4F2F0CDE9086FC63399CB5B659F4C93975819FBD;
defparam prom_inst_11.INIT_RAM_2D = 256'h18C6318C620005B29E8E490E22D25AA28A36B9876E2EE602A5F2EDB6DDC7ED7E;
defparam prom_inst_11.INIT_RAM_2E = 256'h210994D99AAB54CB257D54529400000005554005501505041044451400014413;
defparam prom_inst_11.INIT_RAM_2F = 256'hB8AA156BF9FF3FA1FC3C8113FE7D40E95D3AA176EF9553BE6A0C4621602C2202;
defparam prom_inst_11.INIT_RAM_30 = 256'hFF7291AAC0052814A81241240009FFEFFBF7FFC8A04101E12082802804AFBFFA;
defparam prom_inst_11.INIT_RAM_31 = 256'h24EB49923922807FDFFC01252A955095294A50FEFFEEABFDFDFFFFFEF7FFFFF7;
defparam prom_inst_11.INIT_RAM_32 = 256'hFAABFAAFFFABABBEFE0012090000000E1F90B560EAFAAAFFF0FFEFFE4748172D;
defparam prom_inst_11.INIT_RAM_33 = 256'h255244AB4A97FEFFFFCFFFFFAB0C1FFFA912183FFFF3FFF9112BFFFF3FFF91BE;
defparam prom_inst_11.INIT_RAM_34 = 256'h4EEDD6EDCFFFFFFF6FFFFFFFFFDDBB38670CFF4A975FFB7FDCBF729244890120;
defparam prom_inst_11.INIT_RAM_35 = 256'h2187955540000000000012257DF7EDDDE3311334895F75F2DDAB5FFFD5AB4EEB;
defparam prom_inst_11.INIT_RAM_36 = 256'h00AFD7EFEAAFF7F909280556AB72402BF5F85557F5FFFFFDF9FBFFF20106EB2E;
defparam prom_inst_11.INIT_RAM_37 = 256'hD76BB9FDFBF5FABDDAAA40AEFD4AA54AA55520252975FFB85C2BFFFDC2E1E125;
defparam prom_inst_11.INIT_RAM_38 = 256'h44A529294BC7F291294A420940942EEABFCAA2A945554AA9200000000576BBAE;
defparam prom_inst_11.INIT_RAM_39 = 256'h24A5294A46FFFFFFFC9294A529400011294A52948FFFFFFFFF0494A5294A0A85;
defparam prom_inst_11.INIT_RAM_3A = 256'h4A04A17194929524A5E2A4A4940A12812871A1294252F142502508CA42502502;
defparam prom_inst_11.INIT_RAM_3B = 256'hAAA89294A5294150A82A153D05441281285DF1684210A8052A014BCA92925228;
defparam prom_inst_11.INIT_RAM_3C = 256'hDEAAAAAAAAAAAEAABEAAAAAAAF2AAFFBFFEAAA835555D5555554AB3080050003;
defparam prom_inst_11.INIT_RAM_3D = 256'h55555555555555501985555406615555DDDDC2AAA8082482482485F777DF7757;
defparam prom_inst_11.INIT_RAM_3E = 256'hF0000242840A050287DFFF7777FE8054A54BCA941B94BE22E44440640077400B;
defparam prom_inst_11.INIT_RAM_3F = 256'h003400000000000529004529005A94E3F1F8000200008A12978A052880020000;

pROM prom_inst_12 (
    .DO({prom_inst_12_dout_w[30:0],prom_inst_12_dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_12.READ_MODE = 1'b0;
defparam prom_inst_12.BIT_WIDTH = 1;
defparam prom_inst_12.RESET_MODE = "SYNC";
defparam prom_inst_12.INIT_RAM_00 = 256'hFFFFFFFFFF57A1BDF69CF7DED750C37947407FF1FBF9F9FBFFFF46FFFFFFF901;
defparam prom_inst_12.INIT_RAM_01 = 256'h3715850A3BAC92DB64B6DB24B647C38FF0E4046CF9D9000003F03DC7F00021F6;
defparam prom_inst_12.INIT_RAM_02 = 256'hAF6A3838090ABD97D733333989041A0D200A406833124277D93E2EFB6480CFAF;
defparam prom_inst_12.INIT_RAM_03 = 256'h010BD018C32E2367DD5C7921E34F1BAE342E32822A028A8A800A208A08020A02;
defparam prom_inst_12.INIT_RAM_04 = 256'h606DCDFFD60E6883D83DDDF6C31A316183EF1789CC4CECCE07CEF76672F1B3B9;
defparam prom_inst_12.INIT_RAM_05 = 256'h63F3FFFEB7473E1CBDDF7DFF6FF1DFDED7D47FBA77E61FEF94079C443511B94B;
defparam prom_inst_12.INIT_RAM_06 = 256'hFFCCB14209C5B809FFFEB185C260C0933E1CAE1E79FACCDE7B9F9AC72668C998;
defparam prom_inst_12.INIT_RAM_07 = 256'hF7E664B3C8444CCCF1CDB51CB9845EE615F064F9D1B4736A278C7C088AA2223C;
defparam prom_inst_12.INIT_RAM_08 = 256'h2625BAC00004444E677124850A74C088A844620C5E9C732FFDDD5A3622D44A7D;
defparam prom_inst_12.INIT_RAM_09 = 256'hDA6DD54E0F99986D9A26264D12C4B668989901CD3B6D80248A0B12688E202D9A;
defparam prom_inst_12.INIT_RAM_0A = 256'h989341F090F3F7305D2014FFCDC0672CD1B18668E84B346C6219A3804B346C60;
defparam prom_inst_12.INIT_RAM_0B = 256'hF84BBF7BC9FCBECD3AF8C08104BC7FF73838998F0CB249240899C2810F000897;
defparam prom_inst_12.INIT_RAM_0C = 256'hE7E64F79218099C30C01234FBB1E331CC01330F8B387FCC5FB28E451440DCCDC;
defparam prom_inst_12.INIT_RAM_0D = 256'hE71198F45C738D183F2C27CE787C6831FCBF31841A3201D3D8E78980F8C5E260;
defparam prom_inst_12.INIT_RAM_0E = 256'h910439C44663D8E71A307E584F9CF0F8D063F97E630834640387B1CEE24C7914;
defparam prom_inst_12.INIT_RAM_0F = 256'h241B480F1A13806646000000010EC0CC0B10E206333333311F0030E38FEE24C7;
defparam prom_inst_12.INIT_RAM_10 = 256'h0000182183A54EFB1FD80A050C631ED818A41679880D8106C203C684E011B006;
defparam prom_inst_12.INIT_RAM_11 = 256'h1E301264088133229887CC4E63220090204408FEFFF01BE1F3071F98C6700800;
defparam prom_inst_12.INIT_RAM_12 = 256'h001C6BFF1605BFC8BA4D97103CCC38440DF98C09110E881B0C30C1961B180996;
defparam prom_inst_12.INIT_RAM_13 = 256'h279879365C40F0E11037E63024443A206C4CB0F10093E627665D901E4F309320;
defparam prom_inst_12.INIT_RAM_14 = 256'h64CCCD9345E666B7BF9C8DA4013F9CE2C02198C50BC4AACC857FFFFFFD90B871;
defparam prom_inst_12.INIT_RAM_15 = 256'h6242226667B2ECCE72479CCB638C50B70C4C07E5A79918026659F39F0BC48F26;
defparam prom_inst_12.INIT_RAM_16 = 256'h2ECCE4FD5F56664B2D48444CCCF65966727C91E732DAE35C6285C3FEFFB33259;
defparam prom_inst_12.INIT_RAM_17 = 256'hC06087E043939007004DCE401B782248C064936640BE4BAF332596A42226667B;
defparam prom_inst_12.INIT_RAM_18 = 256'h4ED186C040482F8E70E006048786F9FCF9AFC40A60E10FC0498187FE83000C3F;
defparam prom_inst_12.INIT_RAM_19 = 256'hE6DAFF83317C6B3010312989F0001894F01F16EFBBB332D605503F8F065E3108;
defparam prom_inst_12.INIT_RAM_1A = 256'h02081DEE63423891A1E892683B0283D150880072F188316F8D1796736C7568F3;
defparam prom_inst_12.INIT_RAM_1B = 256'h77F92C924B3273005A16E03F08A2E8A8C482C10000000000C870D7A09000002B;
defparam prom_inst_12.INIT_RAM_1C = 256'hCC2A26D0183217860973FC7DF83E39BFFE0ADE4FC64DA413897315D3B6CAB268;
defparam prom_inst_12.INIT_RAM_1D = 256'h401370C1099269C9C11D811A18E3C09E2726D1204381C0C0621912780E0F7378;
defparam prom_inst_12.INIT_RAM_1E = 256'h01800810FBF8447288CF82452DD451C0737644CEEF82094B6001C44EF10903C8;
defparam prom_inst_12.INIT_RAM_1F = 256'h001B18209CE6E6A5002020A25EEF90E09C4FC1086C1D8A30661883E4F26E2031;
defparam prom_inst_12.INIT_RAM_20 = 256'h284B0F1F438CCD716EB282695190610F0A8F536E60BA402868DC3B618FE80262;
defparam prom_inst_12.INIT_RAM_21 = 256'h5960D93591FF0412090484780802027CCA490A49C6A1A2E56E38602F338F5B6E;
defparam prom_inst_12.INIT_RAM_22 = 256'h57982F305E72BCE57982F305F0270C0486EDE036E52F31A11F25AB1150530800;
defparam prom_inst_12.INIT_RAM_23 = 256'h910E455BC60F79460BF0A395ECE57982F305E72BCE57982F305E72BF93BE46CE;
defparam prom_inst_12.INIT_RAM_24 = 256'hE0CF3C0B2C0CCEB2E7708E0177C91E9E552C76BF4DCBDCCBDF0ECF01F8F8C11C;
defparam prom_inst_12.INIT_RAM_25 = 256'h77850C939F22416CFEF4112B4EA18EDE822533CB4A6C3A1BD27C3694986ED86C;
defparam prom_inst_12.INIT_RAM_26 = 256'h0C30C3041001404063B1013191263224C64919F82409CBDF93EE113C978F3099;
defparam prom_inst_12.INIT_RAM_27 = 256'h8701048121E400348008790C80420870820C41071C61851041810C10C10C3043;
defparam prom_inst_12.INIT_RAM_28 = 256'h00000000000000000000000000000000000000000000000001DFE7D7E687034C;
defparam prom_inst_12.INIT_RAM_29 = 256'h56010AAD1A32555554A9550000000000003FE0606060607FE000000000000000;
defparam prom_inst_12.INIT_RAM_2A = 256'hD5B8254EEAA892A24C1065521688B7875CDCF40000C6018B62EA154DC52DB685;
defparam prom_inst_12.INIT_RAM_2B = 256'h00000050555555555550000000055555555000076C66924836D4DC1362A9B826;
defparam prom_inst_12.INIT_RAM_2C = 256'hCCCDDDDDDCCCCD11111111119888DDCCDDCCCCDDDDCCCDDDDCCCCDDD00055500;
defparam prom_inst_12.INIT_RAM_2D = 256'hCBBBA43FC9BBE4779767CB8FF2EE798BF2777CA3FCDDDCCCCCCCDDDDDDDDDCCC;
defparam prom_inst_12.INIT_RAM_2E = 256'hF237CB9DE49FF2E77927FCB37C9CFF2CDF273FC99FF267FC99FF267FCBBBA43F;
defparam prom_inst_12.INIT_RAM_2F = 256'hCFCE2FAC41F3069349980284000840180333333333330180C0603677CB1FE5CD;
defparam prom_inst_12.INIT_RAM_30 = 256'h00033201FE1FEEF183FDFEFF7FBFDFEEDBBF7EFFDFBF7EFDFBE60D269363F3C5;
defparam prom_inst_12.INIT_RAM_31 = 256'h0000000000000000000001ACB49269249A49749E3FFF003FF3F9E79FCF337400;
defparam prom_inst_12.INIT_RAM_32 = 256'hFFFFF23F9C3FFFFFD5557FFFFFE17FE47FFFC1FF91FFFFFF8000000000000000;
defparam prom_inst_12.INIT_RAM_33 = 256'h2AAE80002878287800001144555551FFFFE411E441E17FFFFE8DFE967FFFFFFF;
defparam prom_inst_12.INIT_RAM_34 = 256'h2AEA9ABA9AAF9ABE1BAA9AAAAAAEFFFFAAAEFAAE9EAEBABAAAAE078687868000;
defparam prom_inst_12.INIT_RAM_35 = 256'h2AAE078A0788114111550000000000000A7802780000000011FFC1E47FE40000;
defparam prom_inst_12.INIT_RAM_36 = 256'hFEBF82A80AAA0AA800001AAFAAAE9D561D561D563AAA9AAA80001AAF9BAA9ABE;
defparam prom_inst_12.INIT_RAM_37 = 256'hF2ABEACBEB32ACACF001F555EAABF555E001EAABEAABAB2B800A00026BFEBFEB;
defparam prom_inst_12.INIT_RAM_38 = 256'h0AAA0AAA00280288000202A8022A02A808020A08000002A86B2BFFFFD5552AAA;
defparam prom_inst_12.INIT_RAM_39 = 256'h1D5600001ABE2AAB8AAA0AAA0AAA00AA0AAA0000020802AA0AAA02A802A80AAA;
defparam prom_inst_12.INIT_RAM_3A = 256'h00005AC6000000002AAA80002AAAEAAAAAAB8001E0000000567EB9E00000AAAE;
defparam prom_inst_12.INIT_RAM_3B = 256'h2AA00000800AFFFF8A020AAA00001E0000000000380607E0786056180795789F;
defparam prom_inst_12.INIT_RAM_3C = 256'h188700000AA80000088AEF528007AAAA8007AD5000006000088AAAAAB377AA00;
defparam prom_inst_12.INIT_RAM_3D = 256'h8001B87FF80079CA80000FFE18A07FFEFFFEE060786180001D6000003D7E0000;
defparam prom_inst_12.INIT_RAM_3E = 256'h80101801008017F801418010080107F8786001FE01E01B80000061FE78007861;
defparam prom_inst_12.INIT_RAM_3F = 256'h010080100801008010080100801008010080100801008017F801008010080100;

pROM prom_inst_13 (
    .DO({prom_inst_13_dout_w[30:0],prom_inst_13_dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_13.READ_MODE = 1'b0;
defparam prom_inst_13.BIT_WIDTH = 1;
defparam prom_inst_13.RESET_MODE = "SYNC";
defparam prom_inst_13.INIT_RAM_00 = 256'h10080100801008010080100801008010080100801008017F8010080100801008;
defparam prom_inst_13.INIT_RAM_01 = 256'h18003F1E3F3F3F1E3F3E061A011E171E2132001E008010080100801008010080;
defparam prom_inst_13.INIT_RAM_02 = 256'hEAAAAEFFFFFFFF800072AB81F80000303103313F0F1F01123F1E3F1E3F3F3F3F;
defparam prom_inst_13.INIT_RAM_03 = 256'hD72CD72AAAAAAA80007F8067E000187FE7FFFF98181E6001E0000000002EAE3A;
defparam prom_inst_13.INIT_RAM_04 = 256'h55554AAAAA8007CB5AAAB52D502AAAD55FEAAAAAABAAAA87FFCBEAAAAACBF72C;
defparam prom_inst_13.INIT_RAM_05 = 256'hFF800801087FFF98181FFE4AAAD2AAD3552AAAAAAAF552EED56F556F52D4AFD5;
defparam prom_inst_13.INIT_RAM_06 = 256'h807FFE7FFF9FFFFF81FFFFFFFFFFE02A002AA00000800ADE005E407FFF80007F;
defparam prom_inst_13.INIT_RAM_07 = 256'h557FFE755500007FFF80004BF801FACAAA9FFFFFFF801800001E0621E020067F;
defparam prom_inst_13.INIT_RAM_08 = 256'h552AAAFFFF80007555000000004AAA8000000007862006780600007FFFFE0075;
defparam prom_inst_13.INIT_RAM_09 = 256'h000780000000009F8660000001F555000680004AAAA0060006200660007FFFD5;
defparam prom_inst_13.INIT_RAM_0A = 256'h000000000000000000000000000000000000000000000000000000000000001E;
defparam prom_inst_13.INIT_RAM_0B = 256'h07FFFFDF840DF800DF800FF800FFFFF800000000000000000000000000000000;
defparam prom_inst_13.INIT_RAM_0C = 256'hC0000FFFFF800000000000000000027FFFFBFF003F6002F0000600C0600C0000;
defparam prom_inst_13.INIT_RAM_0D = 256'h003EDFDFED3C3EDFDFEC4008C7FF8C0000C0000CFDFCD3C3EDFDFEC2008C3FF8;
defparam prom_inst_13.INIT_RAM_0E = 256'hFF0C2AA8C3FF8C2AA8C3FF8C0820C0FE0C0000C0000FFFFFFFFFFC0000CFDFCD;
defparam prom_inst_13.INIT_RAM_0F = 256'h04DF9FCC0000C0000FFFFFFFFFFDFFFEFF9FDFF9FDFF9FDFFFFFC2008C3FF8C1;
defparam prom_inst_13.INIT_RAM_10 = 256'hFDFFFEFF9FDFF9FDFF9FDFFFFFC2008C3FF8DF3FEEAD55FFFFFEAD55FFFFFD09;
defparam prom_inst_13.INIT_RAM_11 = 256'hFFFFF8C03FFFFFFFFFF241101C01E020087A1E87E7F80601007FF0300DFFFFFF;
defparam prom_inst_13.INIT_RAM_12 = 256'h84018FC018F801954319FC49954499FC79884018FC018000180001FFFFF00000;
defparam prom_inst_13.INIT_RAM_13 = 256'h0000000000000FE000000000000000000FFFFF8F801954319FC49954499FC798;
defparam prom_inst_13.INIT_RAM_14 = 256'h4000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_13.INIT_RAM_15 = 256'h0FAAAC000D703C00000000000000040000400000000000000000000000040000;
defparam prom_inst_13.INIT_RAM_16 = 256'hCFAAAFD730000FD7300000FC00C303FFCFC000000FAB0F00C0000FFFF7FD7000;
defparam prom_inst_13.INIT_RAM_17 = 256'hC0000CD5500000D5C00005C0C8FFF000C3FFC0000FD7FF5F00000C000D7FDFD7;
defparam prom_inst_13.INIT_RAM_18 = 256'hF000003AB0000CC0F0000000000003FFCCCD5003FAAD73570000000D5AAD70D5;
defparam prom_inst_13.INIT_RAM_19 = 256'hF00005F5503F003FC0EACD30000003FFC0FC0FBAB00039550A95000C0FEAAFC0;
defparam prom_inst_13.INIT_RAM_1A = 256'hA00000000AAA8AAA8AAAB00003F00FC00D5CC00004440BFFA80803C001211003;
defparam prom_inst_13.INIT_RAM_1B = 256'h0BA303F0000000AAA000000005FD55CC0EB0000005550BFFA8080002A2111EAA;
defparam prom_inst_13.INIT_RAM_1C = 256'h0FFFF000000A20000FC3CFBAFAAABCCD500000000FEB7A57A4F8095F835CF770;
defparam prom_inst_13.INIT_RAM_1D = 256'h7FFFF0FFCF70C0000000000030000D700000033550000FFFF7303F0C0C000F00;
defparam prom_inst_13.INIT_RAM_1E = 256'hC33D70FC0DF5D00FDF3EB73C0FD2C0000387FFD1BFD2CFFFFFFFF387FE47FD55;
defparam prom_inst_13.INIT_RAM_1F = 256'hA0000BCA054213C00CFF0DC0BF0F5F0BC000000000000000000003300C3C0000;
defparam prom_inst_13.INIT_RAM_20 = 256'h03FFC0FF00FFC3FFC3FFC0D550FFF5570FF000000000000000000AAA033C5AAA;
defparam prom_inst_13.INIT_RAM_21 = 256'h00000820000002A7C0000FFF20FF03FFC0FF03FFC030F0000D700E40000013FF;
defparam prom_inst_13.INIT_RAM_22 = 256'h00000000000000000000000000040AAAA000080800000FF00000000000080AA0;
defparam prom_inst_13.INIT_RAM_23 = 256'h0000000000000000200200000000000000000000000000000000000000000000;
defparam prom_inst_13.INIT_RAM_24 = 256'hFFFFC39E67FFFFAAAFFEBFAFFFEEFABE00000000000000000000000000000020;
defparam prom_inst_13.INIT_RAM_25 = 256'h1B5C465888F56C3C1B56C218E5F7DF7F501999B1D63EE5CE6319FF7FFFFF7F6F;
defparam prom_inst_13.INIT_RAM_26 = 256'hD5180ED869EA0EAD86EEF981E29F18C6F44446D5B8DE7394B0DDDD6FDF7E3511;
defparam prom_inst_13.INIT_RAM_27 = 256'hC5C89D5B8B8A36B68EFAB71700003C3E3E0003FFFFECCCC8B8D0DBD61D5B8DDD;
defparam prom_inst_13.INIT_RAM_28 = 256'hF7318C7AC088D0CCC9ADFB96FDCB7EE7DCFD6084206B5F5EF8771C1D6AFDD56E;
defparam prom_inst_13.INIT_RAM_29 = 256'hDF80F9C0D52A2A71BDB7FFDDD1E03FD14EE20810206667002777EE71FFB9E630;
defparam prom_inst_13.INIT_RAM_2A = 256'h3333333333B3311333CF7ABF1FC7FBF00023F0FFDDDDD0097DBD9DCDBF80F9E0;
defparam prom_inst_13.INIT_RAM_2B = 256'hBB9BB0CE8F3AA2BAABECFA153EFDFA6EBB6A520BB592C964BACB2CA09FBC103B;
defparam prom_inst_13.INIT_RAM_2C = 256'h0008123A08F98B84D27A1019DEBE9FA694963D6BCEA272ED34BFBFEE31BBE14F;
defparam prom_inst_13.INIT_RAM_2D = 256'h18C6318C620001B61C6D3F8C23F7E620827E3BE2C65113802C16ED3678003280;
defparam prom_inst_13.INIT_RAM_2E = 256'h405D9861E067983838C599184205555550000005554005501505041044451403;
defparam prom_inst_13.INIT_RAM_2F = 256'hA8AA1FCBF9FF3FE1FC288112AA5540E9773FE176FA9FF2BE4408844240480400;
defparam prom_inst_13.INIT_RAM_30 = 256'h00816F5FFFFAD7EB57EDBEDBFFF00000000000295FBEEE1EDF757FD7FAAFBFFB;
defparam prom_inst_13.INIT_RAM_31 = 256'hDB00B66CC6DD118000008EDAD56A876AD6B5A0FBFEBEFFBC0000000108000008;
defparam prom_inst_13.INIT_RAM_32 = 256'hEAABFFFAAAEFEAAFFA000000FFFFFFF30045000015055500180000000037E8D2;
defparam prom_inst_13.INIT_RAM_33 = 256'hDAADBB54B568000000C0000054F2800056EDE0000030000000000003000010BB;
defparam prom_inst_13.INIT_RAM_34 = 256'h110201020000000000000000002244C798F300B56800000023408D6DBB76FEDF;
defparam prom_inst_13.INIT_RAM_35 = 256'h26798AAABFFFFFFFFFFFE2017DD7422264CEECC8807FFFFD0000000000001100;
defparam prom_inst_13.INIT_RAM_36 = 256'hAA1008000000000116C550A8540DAA840201557FF5FFFFFD51FAFF35FE05FE0A;
defparam prom_inst_13.INIT_RAM_37 = 256'h00000000000801402145A05000B458B458A2C400000A000783C000003C1E62D8;
defparam prom_inst_13.INIT_RAM_38 = 256'h0B5AD2D6B4C00D6AD6B40DF6BF68AEFFEA8AA156BA8AB1562000000000000000;
defparam prom_inst_13.INIT_RAM_39 = 256'h535AD6B5A8000000016D6B5AD6800002D6B5AD6B40000000007B6B5AD6B40000;
defparam prom_inst_13.INIT_RAM_3A = 256'hB5FB45D1836D6ADB5A615B5B6A85ED7ED1518ED69DAD30BDAFDA2C85BDAFDAA2;
defparam prom_inst_13.INIT_RAM_3B = 256'h00016D6B5AD6800001C4E200B89BED7ED15571E0000003FAD5FEB4C56D6DA017;
defparam prom_inst_13.INIT_RAM_3C = 256'h5C00000000000155411554555355500000055542AAAA0AAA2AA83B200002AAA8;
defparam prom_inst_13.INIT_RAM_3D = 256'hAAAAAAAAAAAAAA9FFFEAAAA7FFFAAAA9FFFE6555500000000380057D75DD7DDD;
defparam prom_inst_13.INIT_RAM_3E = 256'h32AAA84D7BF5FAFD05D77F77F7D400000AB0D56015603F317FFFFFFFFFFFFF94;
defparam prom_inst_13.INIT_RAM_3F = 256'h002F00000000000AD6FF8AD655156B5FAFD3FFFCAAAA35ED6BF5FA000000FFFF;

pROM prom_inst_14 (
    .DO({prom_inst_14_dout_w[30:0],prom_inst_14_dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_14.READ_MODE = 1'b0;
defparam prom_inst_14.BIT_WIDTH = 1;
defparam prom_inst_14.RESET_MODE = "SYNC";
defparam prom_inst_14.INIT_RAM_00 = 256'hFFFFFFFFFF77B3BDF6DCF7DEDE50C17947553FF0F9FBFBF9FFFE03FFFFFFF901;
defparam prom_inst_14.INIT_RAM_01 = 256'hB799860E7BEDB6DB6492496DB747E39FE2E108B4A95980000003FC3FB3008132;
defparam prom_inst_14.INIT_RAM_02 = 256'h2F7EF878118AEDB55DB3331B88145A0D209A406837104A32C96B2BAF6480DFE5;
defparam prom_inst_14.INIT_RAM_03 = 256'h051B1111C72C232FFFFE79E7E77F39AC046C32A2800A8A20A80A200822022080;
defparam prom_inst_14.INIT_RAM_04 = 256'h40EDC7FFFE1EEC83D06888ECE73B23C98FEB3699CCCECCCC07ECFFE673F331B8;
defparam prom_inst_14.INIT_RAM_05 = 256'hE3F1FFFEF3633E1CFFFF7FB66DB3BFFEFFFE6DB7E3663FFF9807DC641D9BFBDF;
defparam prom_inst_14.INIT_RAM_06 = 256'hFFE491420CC4F809FFFEF18D8661C1B73E1C8E3E78FFC47E6F0F9FC762384B9C;
defparam prom_inst_14.INIT_RAM_07 = 256'h08266593C044444458CDFF1C9D8E5E763DF0EC7380E633FE239C7C0AA888889C;
defparam prom_inst_14.INIT_RAM_08 = 256'h276DBBC66666666E6361326D1A7EC191A8D4240E5F90FB67FDFFFB322654F582;
defparam prom_inst_14.INIT_RAM_09 = 256'hD0FB554E0F9998E5BB276E5D96E496EC9DB9018D3B6D8024820F12EC9F2025BB;
defparam prom_inst_14.INIT_RAM_0A = 256'h9CB763F081F3ED7C3520247FC5C1472DD93B86ECF84B764EE21BB3C04B764EE0;
defparam prom_inst_14.INIT_RAM_0B = 256'hFC4FBFFF41FCBECD3BB8C18105BC7FFE7C3999DE1D965B6401D9C2810F120897;
defparam prom_inst_14.INIT_RAM_0C = 256'hE3E67FF9218099C30C01234BFF1A7B96C8333878B30FFCCDFBF9E05122089589;
defparam prom_inst_14.INIT_RAM_0D = 256'hA21198E414528718FF2463CE78783871FCBF30943E1201D1D9FF9981FC84E661;
defparam prom_inst_14.INIT_RAM_0E = 256'h80042884466390A50E31FE48C79CF0F070E3F97E61287C240383B3FCA67E7804;
defparam prom_inst_14.INIT_RAM_0F = 256'h6E39DC4E1A13984ECF0494104A0ECCC51B08E104044000040F0020E38FCA67E7;
defparam prom_inst_14.INIT_RAM_10 = 256'hC0BBF8A183A54AFF17FC0A0508E73ED818841ED98B1C938E67138684E613B062;
defparam prom_inst_14.INIT_RAM_11 = 256'h7E7013E4188331679847CCE62120948420C419FBFBF09BF3F3071D90EFF39602;
defparam prom_inst_14.INIT_RAM_12 = 256'h777CEFB717059BC87E7C8530FCEE304C3DF984801104987B8E38C9967B380996;
defparam prom_inst_14.INIT_RAM_13 = 256'h3F8CDB3214C3F0C130F7E61200441261ECECB3F3809FE673725C913E7F19B3E2;
defparam prom_inst_14.INIT_RAM_14 = 256'h64CCCC9644A22212958C50A010BF9C624021B8451B4CABCC8401020FFC906873;
defparam prom_inst_14.INIT_RAM_15 = 256'h22022222229264C6724F8CD9238451B60C5C07E4879008022208B19F0B869F26;
defparam prom_inst_14.INIT_RAM_16 = 256'h264C65C000026659654044444452492632FC93E33648E15C228DA200001332CB;
defparam prom_inst_14.INIT_RAM_17 = 256'hC060876043139047054DCE411378A744C06D9EE6007E5451332CB22022222229;
defparam prom_inst_14.INIT_RAM_18 = 256'h6FC98640404DBF8670E047048786F8DEF9FD840260E10DC0698186DC83008E36;
defparam prom_inst_14.INIT_RAM_19 = 256'hA6DBFB01397C693010733B89F008399DF01F96AD111111B60DF0ED8706DE3100;
defparam prom_inst_14.INIT_RAM_1A = 256'h000C3BF63302714DE0FD926C7B03C1E351A840E9B890397BAD0396F96CFFECD2;
defparam prom_inst_14.INIT_RAM_1B = 256'h77DB6596D93E72805794A07D08E2B9A8C588C02B5EA57B9DC87085203000003E;
defparam prom_inst_14.INIT_RAM_1C = 256'h8E7F6ED8183237865BD3FCFFFC3F3FBFFA1BDEDF4EDDB412925337879FCAF6EC;
defparam prom_inst_14.INIT_RAM_1D = 256'h401020411913F9CFC11D811B1871C4DE636EDBA26703C1E0E03953F80E1FD1F9;
defparam prom_inst_14.INIT_RAM_1E = 256'h01D81D04FFF8663BCEC780060DF041C077F244448E0209CF2001CCCEF08803C8;
defparam prom_inst_14.INIT_RAM_1F = 256'h001B18209CE67666020202035FEF90E09CEDC108461C8310461987E7F3EF403B;
defparam prom_inst_14.INIT_RAM_20 = 256'h00030E3FC69E59D3FEF78E6BF1B0E73F9F9FF75AF86A404879F430E39DA80262;
defparam prom_inst_14.INIT_RAM_21 = 256'h70487DF7BDF606130984C0F03120843E7EC90EC0C6A137E5EE1C206F318B5B6F;
defparam prom_inst_14.INIT_RAM_22 = 256'h97BDAF7B5EF6BDED7B92F725F0771C04A6CDE036C1AFF1A912013F33F0774802;
defparam prom_inst_14.INIT_RAM_23 = 256'h9A0E699FEE4F798E4BF0C725E5C97BDAF7B5EF6BDED7B92F725EE4BF97BE67DC;
defparam prom_inst_14.INIT_RAM_24 = 256'hF25F180A080845E3A7700A0797CB1899316F7CAEDD6BFCEBFFDECF01F9F9871C;
defparam prom_inst_14.INIT_RAM_25 = 256'h338508051FA64044BEFCB12FCFE1889F962597C2CEE41E37F33C659D8839B8DC;
defparam prom_inst_14.INIT_RAM_26 = 256'h2000000000004B4863B01173B32E7665CEF911D8344DCBDFF3FE19BC93C73099;
defparam prom_inst_14.INIT_RAM_27 = 256'h870125C169E80805881A7A0D00C18600618038E0821860820828208208208208;
defparam prom_inst_14.INIT_RAM_28 = 256'h00000000000000000000000000000000000000000000000001F56DFFE687034C;
defparam prom_inst_14.INIT_RAM_29 = 256'h5E080ABD37EA5555542955000000000000000F000F0000002000000000000000;
defparam prom_inst_14.INIT_RAM_2A = 256'h8FB80DCEDE1980001C18EF760D996D835CDCFC0081C4038A73FA1F4F451BEC05;
defparam prom_inst_14.INIT_RAM_2B = 256'h0000005055555555555555555550000000000007D9DDB6C8EDF7B8F1C1EF71E3;
defparam prom_inst_14.INIT_RAM_2C = 256'hCCCDDDDDDDDDDC00000000008888DDCCDDDDDDCCCCCCCDDDDDDDDCCC00000000;
defparam prom_inst_14.INIT_RAM_2D = 256'hDFFFEFFFDFFFEFFFBFFFDFFFF7FFFBFFF7FFFDFFFDCCDDDDDDDDCCCCCCCCCCCC;
defparam prom_inst_14.INIT_RAM_2E = 256'hF7FFDFFFEFFFF7FFFBFFFDFFFDFFFF7FFF7FFFDFFFF7FFFDFFFF7FFFDFFFEFFF;
defparam prom_inst_14.INIT_RAM_2F = 256'h8004600C018307FBFD80028C0008C0180333333333330180C0603FFFDFFFEFFF;
defparam prom_inst_14.INIT_RAM_30 = 256'h000333FE01E7EEFDFBFDFEFF7FBFDFEFDFBF7EFFDFBF7EFDFB060FF7FB20028C;
defparam prom_inst_14.INIT_RAM_31 = 256'h00000000000000000000010C3FFF7FFFDFFFA498351400600201041008373044;
defparam prom_inst_14.INIT_RAM_32 = 256'h7FFF9C3F9C3FFFFF800000007FE57FE4000051FF91FF80000000000000000000;
defparam prom_inst_14.INIT_RAM_33 = 256'h2EAA8000287828780000114400000000000011E451E500007E967E967FFF8000;
defparam prom_inst_14.INIT_RAM_34 = 256'h2AAA9AAA9ABF9ABE1AAA9AAAAEAA80002EAAFEAA9EAAAAAAAAAE078287828000;
defparam prom_inst_14.INIT_RAM_35 = 256'h2AAE07880788114500000000000000000278027800000060000051E400000000;
defparam prom_inst_14.INIT_RAM_36 = 256'hAE9A80000000000000001ABFAEAA9D561D561D562AAA9AAA80001ABF9AAA9ABE;
defparam prom_inst_14.INIT_RAM_37 = 256'hEB2DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000069AE9AE9;
defparam prom_inst_14.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000006AADFFFFD5552AAA;
defparam prom_inst_14.INIT_RAM_39 = 256'hFD57FFFFFABE2EAB800000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_3A = 256'h00005AC600000000200000007FFFFFFFFFFFE001E00060005807E0000000AAAF;
defparam prom_inst_14.INIT_RAM_3B = 256'h2AAA000000AAFFFF8000000000000000000000006001F80067FFDAC600017A07;
defparam prom_inst_14.INIT_RAM_3C = 256'h1A07000002A00000088AEF5500002AAAFFF8554180000000088AAAAAB377A800;
defparam prom_inst_14.INIT_RAM_3D = 256'h800039AF800007CA80000EBE06BFF866F86601FE7861800067FE000067BE0000;
defparam prom_inst_14.INIT_RAM_3E = 256'h0000000000000000000000000000780067FFFE0001F80280000006BE00007861;
defparam prom_inst_14.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_15 (
    .DO({prom_inst_15_dout_w[30:0],prom_inst_15_dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_15.READ_MODE = 1'b0;
defparam prom_inst_15.BIT_WIDTH = 1;
defparam prom_inst_15.RESET_MODE = "SYNC";
defparam prom_inst_15.INIT_RAM_00 = 256'h000000000000000000000000007E000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_02 = 256'hAAAEAA80007FFF8001FFFF800000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_03 = 256'hD72CD72AAAAAAAFFFFFFE066607F807FE7FFFF87E000000000000000002AAE2A;
defparam prom_inst_15.INIT_RAM_04 = 256'h5555552AAAFFFAD4D6D5555541AAAAD2BD2AAAFFFF2AAA87FFAA9AAAAAAA9F2C;
defparam prom_inst_15.INIT_RAM_05 = 256'hFFD50801087FFF8000000052AAAAAAAAD4AAAAAAAACACAFF556F556F5552AAD5;
defparam prom_inst_15.INIT_RAM_06 = 256'hE000007FFFFFFFFFF800007FFFFFF828002AAA000000AADE555E407FFFD5557F;
defparam prom_inst_15.INIT_RAM_07 = 256'h5500007555000000007FFFCAFE0007CAAAFEAA800007FE7FFE01867E00200621;
defparam prom_inst_15.INIT_RAM_08 = 256'h552AAAFFFF80007555000000004AAA80078000006620062006000000007FE01D;
defparam prom_inst_15.INIT_RAM_09 = 256'h000000000000009E18000000007FFF800180007FFFA00600007FFE00007FFFD5;
defparam prom_inst_15.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000400008000000;
defparam prom_inst_15.INIT_RAM_0B = 256'h080000005B6005F6007FF007FF000007FFFF8000040000000002000000000000;
defparam prom_inst_15.INIT_RAM_0C = 256'h000000000000000000003F8FE0080000000400FFC09EFC0FFFF9EF2F0FB3C000;
defparam prom_inst_15.INIT_RAM_0D = 256'h3AC0002000C2C00020000000000000000000000002000C2C0002000000000000;
defparam prom_inst_15.INIT_RAM_0E = 256'h0000155000000015500000000000000000000000000000000000000000002000;
defparam prom_inst_15.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_10 = 256'h00000000000000000000000000000000000000000152AA00000152AA00000000;
defparam prom_inst_15.INIT_RAM_11 = 256'h0000003FC000000800078100000000200802008060180601007FFFFFFFFF8000;
defparam prom_inst_15.INIT_RAM_12 = 256'h000000000000000A800000000A80000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_13 = 256'h00301003010030100301003010030100300000000000A800000000A800000000;
defparam prom_inst_15.INIT_RAM_14 = 256'h007FFC001003010030100301003010030100301003010030100301003FD00301;
defparam prom_inst_15.INIT_RAM_15 = 256'h0FAAA0000FC03000000007FFFE49216492007FFC000000000007FFFE4922E492;
defparam prom_inst_15.INIT_RAM_16 = 256'h0FAAA0FC000000FC00000F00000000000FCFF00000EB003000000FFFF35D3000;
defparam prom_inst_15.INIT_RAM_17 = 256'h0000003D70000CD700000F0038FFF00000000C0005D350F0000007000D35D0FC;
defparam prom_inst_15.INIT_RAM_18 = 256'hC000003AB0000F00C0000000000000000C03500D5AAD735C000000355AAD7CD7;
defparam prom_inst_15.INIT_RAM_19 = 256'hF00005F55000000000EACFC0000000000F0003EAF00009550A9500030F3AAF00;
defparam prom_inst_15.INIT_RAM_1A = 256'h000003F000AA0AA80EAAB0000D5C00000357F00004440AAAA22220FD5020003F;
defparam prom_inst_15.INIT_RAM_1B = 256'h01E1C000000000002000000005FD5F03FEB0000005550AAA8222255552001000;
defparam prom_inst_15.INIT_RAM_1C = 256'h008080000008A0000F0333EACEAABC03500000000FEB7A57A470155140F00770;
defparam prom_inst_15.INIT_RAM_1D = 256'hFFFFF0FFC0FF000000000FFFE0000FC00000000D70000FFFFC0FC003070007C0;
defparam prom_inst_15.INIT_RAM_1E = 256'h303C7F000DD55000F57DBC000FD2C0000387FFD2CFD2CFFFF0000387F387FFFF;
defparam prom_inst_15.INIT_RAM_1F = 256'h000003CA0FF203C003FC0DD6B3FFFAFAC000000000000000000003C00C300000;
defparam prom_inst_15.INIT_RAM_20 = 256'h0000000000000000000000FF70000FD7000000000000000000000555500F0000;
defparam prom_inst_15.INIT_RAM_21 = 256'h000AA2200000000570000FFF2000000000000000000F00000FF00E4000001000;
defparam prom_inst_15.INIT_RAM_22 = 256'h000040000044004000000000000400A000000222200000A00000000000080000;
defparam prom_inst_15.INIT_RAM_23 = 256'h0004000400040040000000000000400400400040000004000004004000044040;
defparam prom_inst_15.INIT_RAM_24 = 256'h6FFFE73446FD5555500055551545141500000000000000000000400400000404;
defparam prom_inst_15.INIT_RAM_25 = 256'h1315EF7CC8FECA0A136CA3D2B5F7DF7FFC9999257088A35EF7BDFFBFDFFF924B;
defparam prom_inst_15.INIT_RAM_26 = 256'hBA87EC91047106D945DDFE001EC40000B44444DB20BF7BDE20BBBB9145362511;
defparam prom_inst_15.INIT_RAM_27 = 256'h8FCC9FB2020B20A0869B6404000003FFC00000000011555F20BA08E20DB28BBB;
defparam prom_inst_15.INIT_RAM_28 = 256'hFF7BDE7E8088D0CCC9A1C390E1C870E11CE056F7BDCADE52F837381C6295F14A;
defparam prom_inst_15.INIT_RAM_29 = 256'hD94495E2D5AB2A51BFFFFFFC91D10C004AE2081020666602256FEF79FFFDE210;
defparam prom_inst_15.INIT_RAM_2A = 256'h333333233112311137DF5AAF3FCF56D0082361FB75555005F92545ED794495E2;
defparam prom_inst_15.INIT_RAM_2B = 256'h92A2A0878D302038025CD2000D9B3658FFFE2303B1D8EC7638E38E20D6DC1003;
defparam prom_inst_15.INIT_RAM_2C = 256'h00001B1E08D98B02D238001015B5836406847BCAC633536B341366E231226043;
defparam prom_inst_15.INIT_RAM_2D = 256'h18C6318C620005241C29128C23450620825A22C0A6599880281CB92430022020;
defparam prom_inst_15.INIT_RAM_2E = 256'h003E603E061FE007C03BE108C605555555555550000005554005501505041043;
defparam prom_inst_15.INIT_RAM_2F = 256'h005400040000154000000000002A80402A000022000000140801008000000000;
defparam prom_inst_15.INIT_RAM_30 = 256'h001290A000052814A812412400080020200000448000000000000000044D4074;
defparam prom_inst_15.INIT_RAM_31 = 256'h24A848922922C848548641252A955095294A5B34C00C53408028140022000000;
defparam prom_inst_15.INIT_RAM_32 = 256'hC00155555507141D000012090000000988000000000000004C24250321080125;
defparam prom_inst_15.INIT_RAM_33 = 256'h255244AA48954A244B6002448904400489120D8912D8912C9128912D8912C931;
defparam prom_inst_15.INIT_RAM_34 = 256'h44894489448912252A4A912A404891202404AA48955529525489520244890120;
defparam prom_inst_15.INIT_RAM_35 = 256'h0004C0000000000000001932EBAEA555300000064C9861820C89448944894489;
defparam prom_inst_15.INIT_RAM_36 = 256'h00A050240028140C8928050281224028140D8002A0AAAAA82801009A01B201B0;
defparam prom_inst_15.INIT_RAM_37 = 256'h000009554A954A954AAA4CAAA54AA54AA5553625295000A0502A800502813125;
defparam prom_inst_15.INIT_RAM_38 = 256'h44A529294A625291294B62094096D554544512A945554AA99000000004000080;
defparam prom_inst_15.INIT_RAM_39 = 256'h24A5294A4494A529489294A529400011294A529484A5294A520494A5294A0A85;
defparam prom_inst_15.INIT_RAM_3A = 256'h4A04B60094929524A53284A494CA12812DA82129425299425025B00A42502530;
defparam prom_inst_15.INIT_RAM_3B = 256'h00009294A5294150A82A1505054412812D88A8884210A80528014A6A12925B28;
defparam prom_inst_15.INIT_RAM_3C = 256'h18AAAAAAAAAAAAAAAAAAAAAAADAAAAAAAAAAAAD9555555555556D40080050001;
defparam prom_inst_15.INIT_RAM_3D = 256'h55555555555555400005555000015554000132AAA80824824826526062206A20;
defparam prom_inst_15.INIT_RAM_3E = 256'h98000322840A0502DB8EA2EA2E228054A54A6A96CA96C0028000000000000008;
defparam prom_inst_15.INIT_RAM_3F = 256'h001B00000000000529004529004A94A05028000200008A12940A052880020000;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_0 (
  .O(dout[0]),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_1_dout[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_1 (
  .O(dout[1]),
  .I0(prom_inst_2_dout[1]),
  .I1(prom_inst_3_dout[1]),
  .S0(dff_q_0)
);
MUX2 mux_inst_2 (
  .O(dout[2]),
  .I0(prom_inst_4_dout[2]),
  .I1(prom_inst_5_dout[2]),
  .S0(dff_q_0)
);
MUX2 mux_inst_3 (
  .O(dout[3]),
  .I0(prom_inst_6_dout[3]),
  .I1(prom_inst_7_dout[3]),
  .S0(dff_q_0)
);
MUX2 mux_inst_4 (
  .O(dout[4]),
  .I0(prom_inst_8_dout[4]),
  .I1(prom_inst_9_dout[4]),
  .S0(dff_q_0)
);
MUX2 mux_inst_5 (
  .O(dout[5]),
  .I0(prom_inst_10_dout[5]),
  .I1(prom_inst_11_dout[5]),
  .S0(dff_q_0)
);
MUX2 mux_inst_6 (
  .O(dout[6]),
  .I0(prom_inst_12_dout[6]),
  .I1(prom_inst_13_dout[6]),
  .S0(dff_q_0)
);
MUX2 mux_inst_7 (
  .O(dout[7]),
  .I0(prom_inst_14_dout[7]),
  .I1(prom_inst_15_dout[7]),
  .S0(dff_q_0)
);
endmodule //cart_prom
